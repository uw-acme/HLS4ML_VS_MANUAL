// Width: 19
// NFRAC: 9
package dense_3_19_9;

localparam logic signed [18:0] weights [32][32] = '{ 
{19'b1111111111111100110, 19'b1111111111100100000, 19'b1111111111100110000, 19'b1111111111110011110, 19'b0000000000010101111, 19'b0000000000000010110, 19'b1111111111111111001, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000001000000, 19'b1111111111011110010, 19'b1111111111111100001, 19'b0000000000110110001, 19'b1111111111110000100, 19'b1111111111000100010, 19'b1111111111111101101, 19'b0000000000000111001, 19'b0000000000011011110, 19'b1111111111101001101, 19'b1111111110111011110, 19'b1111111111111101000, 19'b0000000000000011001, 19'b1111111111100110001, 19'b0000000000000000000, 19'b0000000001000000110, 19'b1111111110100010110, 19'b1111111111110001110, 19'b1111111111100111001, 19'b1111111111110110011, 19'b0000000000011011000, 19'b1111111111110101110}, 
{19'b0000000000101111110, 19'b0000000001101110101, 19'b0000000000011001101, 19'b1111111111010101111, 19'b0000000000001111101, 19'b1111111111101110100, 19'b1111111111111001000, 19'b0000000001000101110, 19'b0000000000000000011, 19'b1111111111111111111, 19'b1111111111111101111, 19'b1111111111011010010, 19'b1111111111110011000, 19'b0000000000100010100, 19'b1111111101111001001, 19'b1111111111100001110, 19'b1111111111111111111, 19'b1111111111111111011, 19'b1111111111111100101, 19'b1111111111110101011, 19'b1111111111101111011, 19'b1111111111101110011, 19'b0000000000000001000, 19'b1111111111111111111, 19'b1111111111111111100, 19'b1111111110111011011, 19'b0000000000000000110, 19'b0000000000011110001, 19'b1111111111111011111, 19'b1111111111010011110, 19'b0000000000000000001, 19'b0000000000000010011}, 
{19'b1111111111000000111, 19'b0000000000001011110, 19'b0000000000000000101, 19'b0000000000010100101, 19'b1111111111010111101, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111001010010, 19'b0000000000100010010, 19'b1111111111101111001, 19'b1111111111101111011, 19'b1111111110100000110, 19'b1111111111101100000, 19'b0000000000100000101, 19'b0000000000010000111, 19'b1111111111111111111, 19'b1111111111111000101, 19'b1111111111111110011, 19'b1111111111001011110, 19'b0000000000000000001, 19'b0000000000000111111, 19'b0000000000000100011, 19'b0000000000001101011, 19'b0000000000111000010, 19'b0000000000000010011, 19'b1111111111001101100, 19'b0000000000110001000, 19'b0000000000000000000, 19'b0000000000001010100, 19'b1111111111111110100, 19'b0000000000000000000, 19'b0000000010010001001}, 
{19'b0000000000110101100, 19'b1111111111111111111, 19'b1111111111110011100, 19'b0000000001010011110, 19'b0000000001001110100, 19'b0000000000000000000, 19'b0000000000000100101, 19'b0000000000110100000, 19'b1111111111100110101, 19'b1111111111111111111, 19'b1111111111001011010, 19'b0000000000000111101, 19'b0000000000010001000, 19'b1111111111010000001, 19'b0000000000000101111, 19'b1111111111110101110, 19'b1111111111111111111, 19'b1111111111101000101, 19'b0000000000000010011, 19'b0000000000000011100, 19'b0000000000000001000, 19'b1111111111111011010, 19'b0000000001001100011, 19'b0000000000101011111, 19'b0000000000101010001, 19'b0000000000011111110, 19'b0000000000101011101, 19'b0000000000000000000, 19'b1111111111111000011, 19'b0000000000111001111, 19'b0000000000011111111, 19'b1111111111110100110}, 
{19'b0000000001000000000, 19'b1111111111111010000, 19'b1111111111010011101, 19'b1111111110011111110, 19'b0000000000111101000, 19'b0000000000000000000, 19'b1111111111001011011, 19'b1111111111011011110, 19'b1111111111111010000, 19'b1111111110011000011, 19'b1111111101110010100, 19'b0000000000111100100, 19'b0000000001010101100, 19'b0000000001000010111, 19'b1111111110110110011, 19'b1111111110011100110, 19'b0000000000000000000, 19'b1111111111101101111, 19'b0000000000011001101, 19'b0000000000010001110, 19'b1111111111100111111, 19'b1111111111111111001, 19'b0000000001011100010, 19'b1111111101010000000, 19'b0000000000001011010, 19'b1111111110101011101, 19'b0000000000001000011, 19'b1111111111100000001, 19'b1111111111011001110, 19'b1111111111111111111, 19'b0000000000001000111, 19'b0000000001001010010}, 
{19'b0000000000000101100, 19'b1111111111111010101, 19'b1111111111011000101, 19'b1111111111011110101, 19'b0000000000101111100, 19'b0000000000000000000, 19'b1111111111011100001, 19'b1111111111101110100, 19'b1111111111001001001, 19'b1111111111110111110, 19'b1111111111111111111, 19'b0000000000010100100, 19'b0000000000000000000, 19'b0000000000101101110, 19'b1111111110111111010, 19'b1111111111101111101, 19'b0000000000001011011, 19'b1111111111011010011, 19'b1111111111100110101, 19'b1111111111111111111, 19'b0000000000000001100, 19'b0000000000100110010, 19'b0000000000111011110, 19'b1111111111111110101, 19'b1111111111111111111, 19'b0000000000110011010, 19'b1111111110111001101, 19'b1111111111111111111, 19'b1111111111100001101, 19'b1111111111111011010, 19'b1111111111111111100, 19'b0000000000000000110}, 
{19'b0000000000001000010, 19'b1111111111010101011, 19'b0000000000001101110, 19'b1111111111111011000, 19'b1111111111111111000, 19'b0000000000010011011, 19'b1111111111110010011, 19'b1111111110101001010, 19'b1111111111111111111, 19'b1111111111100101010, 19'b1111111111000101100, 19'b0000000000111100011, 19'b0000000000000000111, 19'b0000000001010111100, 19'b0000000001101010000, 19'b0000000000000000010, 19'b1111111111111111111, 19'b1111111111010111101, 19'b1111111111111000000, 19'b0000000000100010111, 19'b1111111110011111111, 19'b0000000000010011111, 19'b0000000000101001110, 19'b0000000000000010011, 19'b0000000000010011001, 19'b0000000010011111001, 19'b1111111111001101100, 19'b1111111111110100011, 19'b1111111111100111101, 19'b0000000000111110010, 19'b1111111111111001101, 19'b1111111111101010010}, 
{19'b1111111110110011101, 19'b0000000000000011000, 19'b1111111110101111011, 19'b0000000000110111101, 19'b0000000010000011100, 19'b0000000000001110110, 19'b0000000000000000011, 19'b0000000000000110000, 19'b1111111111111111111, 19'b0000000000010000011, 19'b0000000010100110100, 19'b1111111111111111111, 19'b0000000000110000110, 19'b0000000001001111101, 19'b0000000001100010011, 19'b0000000010000110011, 19'b0000000000000000000, 19'b1111111111000010110, 19'b0000000000101011000, 19'b1111111111111111010, 19'b1111111110101110010, 19'b1111111111100010111, 19'b0000000000000001101, 19'b1111111111110101011, 19'b1111111110111111110, 19'b0000000011110000000, 19'b1111111111100011111, 19'b0000000000000000000, 19'b0000000000000000000, 19'b0000000001110001000, 19'b0000000000001011010, 19'b0000000000110010001}, 
{19'b0000000000110110000, 19'b1111111111111101100, 19'b0000000000000000000, 19'b1111111111111010011, 19'b0000000000001010011, 19'b1111111111111011001, 19'b1111111111111111111, 19'b0000000000010100000, 19'b0000000000011011000, 19'b1111111111011100111, 19'b0000000000010001111, 19'b0000000000010111111, 19'b0000000000000001100, 19'b0000000000101010100, 19'b1111111111100011001, 19'b1111111110011001111, 19'b0000000000000000000, 19'b1111111111111110001, 19'b1111111111111100100, 19'b1111111111000000001, 19'b1111111111111111110, 19'b0000000000000000000, 19'b1111111111100110000, 19'b1111111111111110001, 19'b1111111111110011110, 19'b0000000000010011111, 19'b0000000000101111110, 19'b1111111111110000101, 19'b1111111111111001101, 19'b1111111111111010110, 19'b0000000000000011011, 19'b1111111111001101110}, 
{19'b1111111111101001010, 19'b0000000000110001001, 19'b0000000000000000000, 19'b0000000000000000000, 19'b0000000001100101011, 19'b0000000000101001001, 19'b1111111111111111111, 19'b1111111110111000111, 19'b0000000000001111000, 19'b1111111110100110101, 19'b1111111101001100011, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000110110111, 19'b0000000000001110001, 19'b0000000000000000000, 19'b1111111111010101111, 19'b0000000000000000000, 19'b0000000000000000110, 19'b0000000000000111110, 19'b0000000000011111001, 19'b1111111111111100101, 19'b1111111111010001111, 19'b0000000000000001000, 19'b1111111111111110100, 19'b0000000010001010011, 19'b0000000000101001110, 19'b1111111111111111111, 19'b1111111111110110111, 19'b0000000001010101100, 19'b1111111111111010111, 19'b1111111111110100110}, 
{19'b1111111110111101000, 19'b0000000000010110011, 19'b1111111111111011100, 19'b1111111111111111111, 19'b1111111111100000011, 19'b1111111111001111101, 19'b0000000000000110001, 19'b0000000000010010011, 19'b1111111111111111111, 19'b1111111111101010000, 19'b1111111110110110101, 19'b0000000000011001101, 19'b0000000000100110111, 19'b0000000000000000000, 19'b0000000001101011011, 19'b1111111110111000000, 19'b0000000000001101010, 19'b1111111111001101111, 19'b0000000000100100000, 19'b1111111111111111111, 19'b1111111111111011000, 19'b0000000000001000111, 19'b0000000000001111101, 19'b0000000000000000000, 19'b1111111111000000110, 19'b0000000000000011111, 19'b1111111110111000011, 19'b1111111111111010111, 19'b1111111111111111111, 19'b0000000001010110011, 19'b1111111111100111101, 19'b0000000000000000000}, 
{19'b1111111111111111111, 19'b0000000000001110101, 19'b0000000000000000000, 19'b0000000000110010000, 19'b1111111111110001000, 19'b1111111111111010011, 19'b0000000000000111011, 19'b1111111111111111010, 19'b1111111111111010000, 19'b0000000001010010000, 19'b0000000001011001011, 19'b0000000000000000000, 19'b1111111111010101011, 19'b1111111110100110000, 19'b1111111111111001100, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111110111110, 19'b1111111111000011000, 19'b0000000000110000111, 19'b0000000000000000010, 19'b0000000000101111011, 19'b1111111111111111111, 19'b0000000001000111111, 19'b0000000000001111110, 19'b0000000000100111001, 19'b0000000000111010010, 19'b1111111111111001011, 19'b1111111111001101111, 19'b1111111111000111100, 19'b1111111111111111010, 19'b1111111110101010011}, 
{19'b1111111111100011000, 19'b1111111111111111111, 19'b0000000000001111010, 19'b1111111111001010011, 19'b0000000000001011000, 19'b1111111111111111111, 19'b1111111111100100001, 19'b1111111111111110110, 19'b1111111111101111111, 19'b0000000000000100110, 19'b0000000000001001111, 19'b1111111111110110110, 19'b0000000000000010000, 19'b0000000000011000000, 19'b1111111110101111111, 19'b1111111111100000101, 19'b0000000000011101001, 19'b1111111111101001010, 19'b0000000000000000000, 19'b1111111111111100110, 19'b0000000000011000101, 19'b0000000000000001000, 19'b1111111111111100000, 19'b0000000000000101011, 19'b0000000000100010011, 19'b1111111111110010101, 19'b0000000000000000000, 19'b1111111111000110001, 19'b1111111111100110111, 19'b1111111111111111000, 19'b0000000000010110001, 19'b0000000000000000000}, 
{19'b1111111110111101011, 19'b0000000000110101110, 19'b1111111111111111111, 19'b1111111111111111001, 19'b1111111111111110110, 19'b0000000000010110011, 19'b1111111111111111111, 19'b0000000001100010110, 19'b1111111111111110000, 19'b1111111111111111111, 19'b0000000000011010010, 19'b0000000000000101001, 19'b0000000000000000110, 19'b0000000000000000000, 19'b0000000000001111100, 19'b0000000000101010010, 19'b0000000000010110110, 19'b0000000000010101010, 19'b1111111111111110111, 19'b0000000000100111010, 19'b0000000000001100111, 19'b0000000000000101001, 19'b1111111111111110111, 19'b0000000000100000100, 19'b1111111111110011010, 19'b1111111111010100100, 19'b1111111111110100001, 19'b1111111111111111111, 19'b0000000000001101000, 19'b0000000000000011110, 19'b0000000000011001000, 19'b0000000000111101010}, 
{19'b1111111111111101100, 19'b1111111111001110001, 19'b0000000000000110100, 19'b1111111111111111111, 19'b0000000001110101010, 19'b1111111111100101011, 19'b1111111110110110110, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111111100101, 19'b0000000000000110001, 19'b0000000000110111111, 19'b0000000000101001001, 19'b0000000000000001010, 19'b0000000000000100010, 19'b1111111111101001101, 19'b0000000000000100010, 19'b1111111111111011001, 19'b0000000000000000000, 19'b0000000000001001101, 19'b1111111111111011001, 19'b0000000000000010011, 19'b0000000000100010000, 19'b0000000000000100101, 19'b1111111111111110011, 19'b1111111111001011001, 19'b0000000000011010000, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111110010011, 19'b1111111111111101010, 19'b1111111111110111111}, 
{19'b0000000000000000111, 19'b1111111111110111111, 19'b1111111111101111110, 19'b1111111111100100000, 19'b1111111110111010000, 19'b0000000001001110000, 19'b0000000000000000000, 19'b0000000000010101100, 19'b0000000000100100101, 19'b0000000000000001101, 19'b1111111111111011101, 19'b0000000000111100111, 19'b0000000000011100101, 19'b1111111111010001001, 19'b1111111111101011001, 19'b1111111111111010101, 19'b1111111111001101000, 19'b1111111111111101110, 19'b0000000000000000000, 19'b1111111111111111011, 19'b0000000000010011111, 19'b1111111111101110011, 19'b0000000000000000000, 19'b0000000000001001110, 19'b1111111111111111111, 19'b1111111111010100010, 19'b0000000000010100000, 19'b0000000000000000000, 19'b0000000000000101101, 19'b0000000000000001011, 19'b1111111111010111100, 19'b0000000000000010101}, 
{19'b1111111111100110111, 19'b1111111111101011110, 19'b0000000000001001110, 19'b1111111111110000000, 19'b1111111111110100100, 19'b0000000000001110110, 19'b1111111111111111010, 19'b0000000000000100011, 19'b0000000000010000110, 19'b1111111111111111111, 19'b0000000000001111110, 19'b1111111111101111101, 19'b1111111111111110110, 19'b1111111111111111111, 19'b0000000000001101001, 19'b1111111111111111111, 19'b0000000000111110100, 19'b1111111111111101110, 19'b0000000000011111110, 19'b1111111111101010010, 19'b0000000000010100010, 19'b0000000000001000000, 19'b0000000000001010110, 19'b0000000000000100101, 19'b1111111111110101100, 19'b1111111111011100010, 19'b1111111111011110110, 19'b0000000000001101110, 19'b1111111111110101010, 19'b0000000000000000000, 19'b1111111111111100011, 19'b0000000000011101101}, 
{19'b1111111111111111111, 19'b1111111111001100001, 19'b1111111111001101001, 19'b1111111111111111111, 19'b0000000001010000110, 19'b1111111111110100011, 19'b0000000000000000000, 19'b0000000000111101110, 19'b1111111111101101000, 19'b0000000000000000000, 19'b1111111111001010100, 19'b1111111111000001010, 19'b0000000000111001011, 19'b0000000000010011010, 19'b1111111111110000011, 19'b1111111111011100111, 19'b0000000000010110000, 19'b0000000000000000000, 19'b1111111111100001100, 19'b0000000000000011011, 19'b0000000000001000111, 19'b1111111111110100101, 19'b0000000000100100010, 19'b1111111110000010100, 19'b0000000000000101001, 19'b0000000000011110100, 19'b1111111111111010101, 19'b0000000000000001111, 19'b1111111111100010001, 19'b1111111111111111111, 19'b1111111111100110010, 19'b1111111111111100111}, 
{19'b0000000000011011001, 19'b0000000000101100001, 19'b0000000001000110011, 19'b1111111111100101110, 19'b0000000000110101010, 19'b0000000000100111001, 19'b0000000000000000000, 19'b0000000000111010010, 19'b0000000000101101101, 19'b1111111111110010010, 19'b0000000001011001110, 19'b1111111111010011010, 19'b0000000001001111100, 19'b0000000000111001001, 19'b1111111101110110101, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000000000101, 19'b0000000000100001010, 19'b1111111110111111100, 19'b0000000000011100010, 19'b1111111111100100110, 19'b1111111111000001001, 19'b1111111111101011111, 19'b0000000000101010001, 19'b1111111110101011100, 19'b1111111111010101110, 19'b1111111111111010101, 19'b1111111111111111111, 19'b1111111110110111110, 19'b0000000000110010100, 19'b0000000000000000000}, 
{19'b1111111111111001101, 19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111010011000, 19'b0000000000000001001, 19'b0000000000000001000, 19'b1111111111111110000, 19'b1111111111111100111, 19'b1111111111111010000, 19'b0000000000010001110, 19'b1111111111111111111, 19'b0000000000001010100, 19'b1111111111010100001, 19'b0000000000001101101, 19'b1111111111111111111, 19'b0000000000010010000, 19'b0000000000111001010, 19'b1111111111010010110, 19'b0000000000000110101, 19'b1111111111110011010, 19'b0000000000010000011, 19'b0000000000011000010, 19'b1111111111110101000, 19'b1111111111011111110, 19'b0000000000000010101, 19'b0000000001101010001, 19'b1111111111111100111, 19'b1111111111111110000, 19'b0000000000101001100, 19'b0000000000000000000, 19'b0000000001101110010}, 
{19'b1111111110111101001, 19'b0000000000000100101, 19'b1111111111100100010, 19'b0000000000110001000, 19'b0000000000001110000, 19'b1111111111111011111, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111011001001, 19'b1111111111111011110, 19'b0000000000000000000, 19'b1111111110111000111, 19'b0000000000000001100, 19'b1111111111111010111, 19'b1111111111111111101, 19'b1111111111111111111, 19'b1111111111110001000, 19'b0000000000000000101, 19'b0000000000000000011, 19'b0000000000010100010, 19'b0000000000000010001, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111111110111, 19'b0000000000000000000, 19'b0000000000000010010, 19'b0000000001001010011, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111111010110, 19'b0000000000010110011, 19'b1111111111111100101}, 
{19'b1111111111111111110, 19'b1111111111101100101, 19'b0000000000011010001, 19'b0000000000000101000, 19'b1111111111010000011, 19'b0000000000000000000, 19'b0000000000100100100, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111110011011, 19'b0000000000001110101, 19'b0000000000000010011, 19'b0000000000101001011, 19'b1111111110111001110, 19'b1111111111110011111, 19'b1111111111111101110, 19'b0000000000011011101, 19'b1111111111001110110, 19'b0000000000000010101, 19'b1111111110011111011, 19'b1111111111111101100, 19'b1111111111110000110, 19'b1111111111111010110, 19'b0000000000100101110, 19'b1111111111110110011, 19'b1111111111011100000, 19'b0000000000001011100, 19'b0000000000000000000, 19'b0000000000110010101, 19'b0000000001000010111, 19'b1111111111010110000, 19'b1111111111000110100}, 
{19'b0000000000001000101, 19'b0000000000000011010, 19'b1111111111001010111, 19'b1111111111111000101, 19'b1111111111111111111, 19'b0000000000000000010, 19'b0000000000001101100, 19'b0000000000110100101, 19'b0000000000000000000, 19'b0000000000000010100, 19'b0000000000001000111, 19'b1111111110111010111, 19'b1111111111110111011, 19'b1111111110110010101, 19'b0000000000111101100, 19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111110101101111, 19'b1111111111111111111, 19'b1111111111110110011, 19'b1111111111111101010, 19'b0000000000000000000, 19'b0000000000000111111, 19'b1111111111101100110, 19'b0000000000000110110, 19'b0000000000110100100, 19'b0000000000110110100, 19'b0000000000110001111, 19'b0000000000100111011, 19'b0000000000000000000, 19'b0000000000001110100, 19'b0000000001100100010}, 
{19'b1111111111111100110, 19'b1111111111100001100, 19'b0000000000110001110, 19'b1111111111110010110, 19'b0000000000001000111, 19'b0000000000010101011, 19'b1111111111111111111, 19'b1111111111011011010, 19'b1111111111110101000, 19'b1111111110110011000, 19'b0000000000111001010, 19'b0000000000000000011, 19'b0000000000110101101, 19'b0000000001010101110, 19'b1111111111110001000, 19'b1111111110010000100, 19'b1111111111110010101, 19'b0000000000111100001, 19'b1111111111011011110, 19'b1111111111100101010, 19'b0000000000000111100, 19'b0000000000000000001, 19'b1111111110111010001, 19'b1111111111100111100, 19'b1111111111111010111, 19'b1111111111110000011, 19'b0000000000001110010, 19'b0000000001011010000, 19'b0000000000011111011, 19'b1111111111111111111, 19'b0000000000001010010, 19'b0000000000000011100}, 
{19'b0000000000000101011, 19'b0000000000111010000, 19'b0000000000000000000, 19'b0000000000100101110, 19'b0000000001101010011, 19'b1111111111101010001, 19'b1111111111111111111, 19'b1111111111111010010, 19'b0000000000100101100, 19'b1111111111100111011, 19'b1111111111111111110, 19'b0000000000101010101, 19'b0000000000000001000, 19'b0000000000000011100, 19'b1111111100111100100, 19'b1111111111110101110, 19'b0000000000000000000, 19'b0000000000011001101, 19'b1111111111111111100, 19'b0000000000100110001, 19'b1111111111111111111, 19'b1111111111101001111, 19'b1111111110111000000, 19'b0000000000010000101, 19'b0000000000100100100, 19'b1111111101110010000, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000001000101101, 19'b1111111110011001011, 19'b0000000000000000001, 19'b1111111111111111001}, 
{19'b0000000000000001001, 19'b1111111111010100100, 19'b0000000000000110111, 19'b1111111111111110000, 19'b0000000000000110101, 19'b0000000001000011101, 19'b1111111110100011001, 19'b0000000000000100011, 19'b0000000000110110001, 19'b1111111111010100110, 19'b1111111111111101000, 19'b0000000000000110010, 19'b1111111111111110110, 19'b0000000000010110111, 19'b0000000000001101101, 19'b1111111111111101110, 19'b0000000000001000100, 19'b0000000000000000000, 19'b0000000000000010110, 19'b0000000000110000100, 19'b1111111111111100011, 19'b1111111111000010000, 19'b1111111110110010100, 19'b1111111111100111001, 19'b1111111110110100011, 19'b0000000000011010101, 19'b0000000001001111110, 19'b0000000000101111001, 19'b1111111111111110101, 19'b1111111111010000010, 19'b1111111111011000001, 19'b0000000000000111101}, 
{19'b0000000000000110101, 19'b1111111111000010110, 19'b1111111111111101110, 19'b0000000000010011010, 19'b1111111111000010110, 19'b0000000000010101101, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000100001110, 19'b1111111111111101110, 19'b0000000000000001001, 19'b0000000000000000000, 19'b0000000000010000010, 19'b1111111111111101110, 19'b0000000000000000010, 19'b1111111111111111111, 19'b1111111111010110110, 19'b1111111110111111010, 19'b1111111111111111111, 19'b1111111110111011101, 19'b1111111111011001011, 19'b1111111111010000011, 19'b0000000001110001111, 19'b0000000000000010010, 19'b1111111111111010000, 19'b0000000000101000100, 19'b0000000001110010111, 19'b0000000000110010100, 19'b1111111101111000010, 19'b1111111111101000010}, 
{19'b0000000000110000000, 19'b1111111111111111111, 19'b0000000000100000001, 19'b1111111111111101011, 19'b0000000000111101111, 19'b1111111111101101101, 19'b0000000000001001000, 19'b0000000000110101100, 19'b0000000000100010010, 19'b1111111110111101001, 19'b1111111111111000000, 19'b0000000000001111101, 19'b0000000000001000110, 19'b1111111111111110001, 19'b0000000000001010110, 19'b0000000000000000000, 19'b0000000000101110011, 19'b0000000000000100011, 19'b0000000000101111111, 19'b1111111111110111100, 19'b1111111111101111101, 19'b1111111111110110011, 19'b1111111111111111111, 19'b0000000000100110101, 19'b1111111111100110000, 19'b1111111111111111001, 19'b0000000000000000000, 19'b0000000000000000000, 19'b0000000000000000000, 19'b0000000000100101011, 19'b1111111111010110111, 19'b1111111111111101000}, 
{19'b1111111111111111111, 19'b1111111111111100000, 19'b1111111111000100011, 19'b0000000000100100011, 19'b0000000000011100100, 19'b1111111111110001111, 19'b1111111111111111111, 19'b1111111111100010111, 19'b0000000000000000110, 19'b1111111111111111111, 19'b1111111111011001011, 19'b1111111111100000011, 19'b0000000000111101010, 19'b0000000000000000000, 19'b1111111111101111101, 19'b1111111111111111111, 19'b0000000000011011011, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111100100010, 19'b0000000000101000011, 19'b0000000000000000000, 19'b0000000000010011111, 19'b1111111111111100010, 19'b0000000000010100000, 19'b0000000000000000010, 19'b0000000000000000000, 19'b0000000000011110110, 19'b1111111111100111011, 19'b1111111111111010000, 19'b0000000000010100100, 19'b1111111111110010011}, 
{19'b1111111111111101110, 19'b1111111111011000100, 19'b0000000001001100000, 19'b1111111111110111101, 19'b0000000000011001001, 19'b1111111111011011011, 19'b0000000000000000000, 19'b0000000000000100011, 19'b1111111111000010101, 19'b1111111111111110010, 19'b1111111111110000001, 19'b0000000000000111011, 19'b1111111111010110000, 19'b0000000000010001101, 19'b0000000000011001111, 19'b0000000000001110000, 19'b0000000000001010111, 19'b1111111111111011001, 19'b1111111110100101010, 19'b1111111111111110010, 19'b1111111111111000101, 19'b0000000000010001111, 19'b1111111111110001110, 19'b1111111111111111111, 19'b0000000000011001010, 19'b1111111111111010001, 19'b1111111111111110001, 19'b0000000000110001110, 19'b1111111111001101000, 19'b1111111111011010001, 19'b0000000000101100111, 19'b0000000000000100100}, 
{19'b0000000000110111001, 19'b0000000000011001110, 19'b0000000000000000000, 19'b1111111111101011101, 19'b1111111111110101111, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111110111001, 19'b1111111111110000000, 19'b1111111111110000110, 19'b0000000000000000000, 19'b0000000000010100010, 19'b0000000000000000110, 19'b0000000000000110110, 19'b1111111111111010010, 19'b0000000000000000101, 19'b1111111111101100010, 19'b0000000000000000000, 19'b1111111111111101101, 19'b1111111111111111111, 19'b0000000000000000010, 19'b0000000000000111100, 19'b0000000000001100011, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111110110001110, 19'b1111111111100110011, 19'b0000000000000000110, 19'b0000000000000010100, 19'b0000000000000000001, 19'b1111111111101001010, 19'b0000000000000010101}, 
{19'b0000000000011000000, 19'b1111111101111010010, 19'b1111111111111111111, 19'b1111111111110110010, 19'b1111111111100010001, 19'b1111111111111110110, 19'b0000000000000000000, 19'b0000000001000110000, 19'b1111111111111010011, 19'b1111111111111101001, 19'b0000000000001010100, 19'b1111111110101011011, 19'b0000000000000011000, 19'b1111111111000111111, 19'b0000000001011100011, 19'b1111111111111001010, 19'b1111111111100011000, 19'b1111111110111001111, 19'b1111111111111110101, 19'b1111111110100101011, 19'b1111111110011000010, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000000000000, 19'b0000000000011111001, 19'b1111111111111110001, 19'b1111111111011001110, 19'b1111111111110110101, 19'b1111111111111101000, 19'b0000000000000000000, 19'b1111111111111011111, 19'b1111111110100110011}
};

localparam logic signed [18:0] bias [32] = '{
19'b0000000000100001110,  // 0.5280959606170654
19'b0000000000110101110,  // 0.8414360880851746
19'b0000000000011001011,  // 0.397830605506897
19'b0000000000011010010,  // 0.4105983078479767
19'b1111111100010101111,  // -3.657735586166382
19'b1111111111000110100,  // -0.8977976441383362
19'b0000000001101101001,  // 1.7051936388015747
19'b1111111110101110010,  // -1.2765135765075684
19'b1111111111011010101,  // -0.5837795734405518
19'b0000000010101100110,  // 2.699671983718872
19'b0000000000001101111,  // 0.2170683741569519
19'b0000000000111000011,  // 0.8814588785171509
19'b1111111101010111011,  // -2.634300947189331
19'b1111111110000111110,  // -1.877297282218933
19'b0000000001101010011,  // 1.6625694036483765
19'b0000000010101111101,  // 2.7459704875946045
19'b1111111111100001011,  // -0.47838035225868225
19'b0000000001101100101,  // 1.6984987258911133
19'b0000000000110110101,  // 0.8548859357833862
19'b0000000001000000010,  // 1.0045719146728516
19'b0000000001011010110,  // 1.4197649955749512
19'b0000000000110101010,  // 0.832463800907135
19'b0000000000100010110,  // 0.5434179306030273
19'b0000000000111011010,  // 0.9277304410934448
19'b1111111111101010000,  // -0.3426123857498169
19'b1111111111011100001,  // -0.5587119460105896
19'b1111111111011000010,  // -0.6208624839782715
19'b1111111110101110000,  // -1.2802538871765137
19'b0000000000000011110,  // 0.05940237268805504
19'b1111111111001011011,  // -0.8213341236114502
19'b0000000000111000001,  // 0.8783953189849854
19'b1111111111000011001   // -0.949700653553009
};
endpackage