// Width: 24
// NFRAC: 12
package dense_1_24_12;

localparam logic signed [23:0] weights [16][64] = '{ 
{24'b000000000000010000010100, 24'b111111111111010110010010, 24'b111111111111110100011011, 24'b111111111111110001100000, 24'b111111111111100110000101, 24'b000000000000000111000100, 24'b111111111110111101101000, 24'b000000000000000000000000, 24'b000000000000000011101101, 24'b000000000000010000110111, 24'b000000000000000000001100, 24'b111111111111100110000110, 24'b111111111111111111111011, 24'b000000000000001101011000, 24'b000000000000000010001001, 24'b111111111111101111010000, 24'b000000000000001110111001, 24'b000000000000000011110000, 24'b000000000000000000000000, 24'b111111111111111111111111, 24'b000000000000011000000111, 24'b111111111111101010110010, 24'b111111111111111110100101, 24'b000000000000011110010000, 24'b111111111111101011011011, 24'b111111111111010100010100, 24'b111111111111101110010111, 24'b111111111111110011100000, 24'b111111111111111001010011, 24'b111111111111111111111000, 24'b000000000000000010011010, 24'b000000000000001111101101, 24'b000000000000001100100001, 24'b111111111111111111001010, 24'b000000000000000000000000, 24'b000000000000010011111011, 24'b111111111111111110110110, 24'b111111111111101111111011, 24'b000000000000000001101111, 24'b000000000000001100010100, 24'b111111111111111111001110, 24'b000000000000010001100111, 24'b111111111111101110111100, 24'b000000000000111011011100, 24'b111111111111111111111011, 24'b000000000000011100111101, 24'b000000000000000000000000, 24'b000000000000001011110011, 24'b000000000000001100100011, 24'b111111111111111110011111, 24'b000000000000000000000000, 24'b000000000000001010010001, 24'b000000000000001101110100, 24'b000000000000000100111110, 24'b111111111111111000100111, 24'b111111111111101100001000, 24'b000000000000100010010101, 24'b111111111111100000000001, 24'b000000000000011101111011, 24'b111111111111101001010100, 24'b000000000000110010110000, 24'b111111111111111111100001, 24'b000000000000000000101110, 24'b000000000000000101001100}, 
{24'b000000000000000000001011, 24'b111111111111101011011110, 24'b111111111111110111100001, 24'b111111111111101110000110, 24'b111111111111101011101011, 24'b000000000000000110110100, 24'b111111111111001111101101, 24'b111111111111111111110110, 24'b111111111111110001011101, 24'b000000000000001011000010, 24'b000000000000000000011011, 24'b111111111111111010011111, 24'b000000000000001100100111, 24'b000000000000000000000000, 24'b111111111111111111111111, 24'b000000000000001101010010, 24'b111111111111111111100111, 24'b000000000000000000000001, 24'b111111111111110100010101, 24'b111111111111101111111111, 24'b000000000000011100010011, 24'b111111111111111010110100, 24'b000000000000000011000100, 24'b000000000000101100101110, 24'b000000000000010000011110, 24'b111111111111110001010000, 24'b111111111111110001001110, 24'b111111111111111111111110, 24'b111111111111111001100000, 24'b111111111111100110000011, 24'b111111111111111100001010, 24'b000000000000011101000111, 24'b000000000000010001110101, 24'b000000000000100011001101, 24'b000000000000101000010000, 24'b000000000000000011001110, 24'b111111111111111000011011, 24'b111111111111100100001110, 24'b000000000000000011101000, 24'b000000000000001100000101, 24'b000000000000000001011101, 24'b000000000000001101001101, 24'b111111111111110010011001, 24'b000000000000010000001000, 24'b000000000000001011000001, 24'b000000000000000011001100, 24'b111111111111101010001111, 24'b000000000000000101000101, 24'b000000000000010000101011, 24'b000000000000000001111010, 24'b000000000000000001100101, 24'b000000000001001010000100, 24'b111111111111111011001101, 24'b111111111111111001101110, 24'b111111111111111100100001, 24'b111111111111111111100000, 24'b000000000000010000011100, 24'b111111111111101000010100, 24'b000000000000111111000011, 24'b000000000000000000010011, 24'b000000000000100001010100, 24'b000000000000001111010111, 24'b000000000000110100101001, 24'b000000000000001001000001}, 
{24'b111111111111111111100000, 24'b000000000000000000000000, 24'b111111111111111010101011, 24'b111111111111110100101111, 24'b111111111111110100001011, 24'b000000000000000010101011, 24'b000000000001011110110001, 24'b111111111111111111111111, 24'b111111111110101110111110, 24'b111111111111111111111111, 24'b111111111111111111111000, 24'b111111111111111110110110, 24'b111111111111110001011100, 24'b000000000000000000000101, 24'b111111111111111111011001, 24'b000000000000001010110000, 24'b000000000000111001111100, 24'b111111111111111111111111, 24'b000000000000000100100111, 24'b000000000000000000000001, 24'b000000000000011010011000, 24'b111111111111010001110101, 24'b000000000000100100111101, 24'b111111111111010010010100, 24'b000000000000111100101101, 24'b111111111111101001110101, 24'b111111111111110000010101, 24'b111111111111010010000100, 24'b000000000001010001100000, 24'b000000000000010001101001, 24'b000000000000000000101110, 24'b000000000000100001001000, 24'b000000000001000001010011, 24'b111111111110110011100001, 24'b111111111111111001111000, 24'b000000000000000010000010, 24'b111111111111110001001101, 24'b000000000000111001011010, 24'b111111111111111101011110, 24'b000000000000010100000010, 24'b000000000000010101010100, 24'b000000000000010111101010, 24'b111111111111111111111111, 24'b111111111111111111111111, 24'b111111111111111110111001, 24'b000000000000001010000011, 24'b111111111111101110000110, 24'b111111111111110101000110, 24'b111111111111111110111000, 24'b000000000000011001001011, 24'b111111111111110100101111, 24'b000000000000001001100111, 24'b111111111111111111111110, 24'b000000000000001000100101, 24'b111111111111110100110001, 24'b111111111111111111111111, 24'b111111111111101100010001, 24'b111111111111010101001001, 24'b111111111111111111110111, 24'b000000000000000000000000, 24'b000000000001100010101111, 24'b000000000000000000110101, 24'b111111111111111111110101, 24'b111111111111101100001100}, 
{24'b111111111111100010101011, 24'b111111111111101000011010, 24'b111111111111010011101010, 24'b000000000000010011101110, 24'b111111111111101011110010, 24'b111111111110101001110101, 24'b111111111111111000101010, 24'b111111111111101100010010, 24'b000000000000001110010101, 24'b111111111111111111111111, 24'b000000000001010000111111, 24'b111111111111111001001111, 24'b111111111111001101111011, 24'b000000000000100101000100, 24'b000000000000000001100111, 24'b111111111111111111111001, 24'b111111111111100011100110, 24'b111111111111111111111111, 24'b000000000000000000000000, 24'b111111111111110001100001, 24'b111111111110110110010101, 24'b111111111111111000110110, 24'b111111111111010011010011, 24'b000000000000001100101100, 24'b111111111111100111001111, 24'b111111111111000101000101, 24'b000000000000010100000001, 24'b000000000000101111001001, 24'b000000000001010010111001, 24'b111111111111100010100100, 24'b111111111111011010101101, 24'b000000000000000100101110, 24'b000000000000100000000000, 24'b111111111111001010001010, 24'b111111111111101011111000, 24'b000000000000000000000000, 24'b111111111111010001100010, 24'b000000000000001111100001, 24'b111111111111100011110001, 24'b000000000000000111101000, 24'b000000000000011101010110, 24'b000000000000001010000010, 24'b000000000000000000000000, 24'b000000000000000001010011, 24'b000000000000100011010111, 24'b111111111111110011001101, 24'b111111111111111111111111, 24'b111111111111101001111111, 24'b111111111111111111111111, 24'b111111111111111001110011, 24'b111111111111011000100111, 24'b000000000000000101100011, 24'b111111111111111111111111, 24'b000000000000001101111101, 24'b000000000000010100001011, 24'b000000000000101001011010, 24'b111111111111000010000100, 24'b111111111111000100100011, 24'b111111111111010010110111, 24'b000000000000110111011100, 24'b000000000001101111111100, 24'b111111111111000110011011, 24'b111111111111111100100010, 24'b000000000000011011110010}, 
{24'b000000000000010101111001, 24'b111111111111011000011010, 24'b111111111111101111011001, 24'b111111111111111111111111, 24'b111111111111110110001001, 24'b000000000000010101110001, 24'b000000000000001100001000, 24'b111111111111111111111111, 24'b111111111111011001110001, 24'b111111111111110000100001, 24'b111111111111101000011001, 24'b000000000000000011011000, 24'b000000000000000000000101, 24'b000000000000000000000000, 24'b111111111111111101011010, 24'b000000000000010110111000, 24'b000000000000001000100011, 24'b111111111111100110110110, 24'b000000000000000001111101, 24'b000000000000000000110111, 24'b000000000000001101011100, 24'b111111111111111000011100, 24'b000000000000000100110000, 24'b111111111111111110110001, 24'b000000000001000100001101, 24'b111111111111110100000100, 24'b111111111111101110000000, 24'b111111111111100110001010, 24'b000000000000000000000000, 24'b000000000000001010100010, 24'b000000000000000111011100, 24'b000000000000010001100000, 24'b111111111111111111001101, 24'b000000000000000100101111, 24'b000000000000001000010111, 24'b111111111111111111111111, 24'b000000000000000000011001, 24'b000000000000111000011010, 24'b111111111111101101100000, 24'b111111111111111011000110, 24'b000000000000011011101110, 24'b000000000000001111111011, 24'b111111111111100000101101, 24'b000000000000000000011000, 24'b111111111110111011101000, 24'b111111111111111111111111, 24'b111111111111111000001010, 24'b000000000000000000110000, 24'b111111111111111111111111, 24'b111111111111111110011111, 24'b111111111111111111111111, 24'b000000000000001100000010, 24'b111111111111111111101011, 24'b000000000000010100010101, 24'b111111111111110011110001, 24'b111111111111010000111100, 24'b111111111111100010001001, 24'b111111111111011111011001, 24'b111111111111011000101101, 24'b000000000000101111110011, 24'b000000000001010111111010, 24'b000000000000110010101111, 24'b000000000000000111110110, 24'b111111111111111111111111}, 
{24'b111111111111100011011110, 24'b111111111111010111101001, 24'b000000000000000000000000, 24'b000000000000010011101010, 24'b000000000000010010010000, 24'b111111111111110010011011, 24'b000000000000100101010000, 24'b111111111111111111111111, 24'b000000000000001111100110, 24'b111111111111111111111111, 24'b111111111111111111011001, 24'b111111111111111011010110, 24'b111111111111110100101101, 24'b000000000000100101000000, 24'b111111111111111010010010, 24'b000000000000000000000000, 24'b111111111111011000000000, 24'b111111111111101001010100, 24'b000000000000000000000000, 24'b111111111111111111111111, 24'b111111111111111100111101, 24'b111111111111101011111010, 24'b111111111111101011100110, 24'b000000000000011101110010, 24'b111111111111101011101001, 24'b111111111111111111111100, 24'b000000000000010000011001, 24'b111111111111111011010100, 24'b111111111111000100010011, 24'b111111111111111111111111, 24'b111111111111111011101110, 24'b111111111111111111010101, 24'b111111111111111111010000, 24'b000000000000000010100111, 24'b000000000000001000011100, 24'b000000000000010110001000, 24'b000000000000000000110111, 24'b111111111111111001101110, 24'b111111111111101111001100, 24'b111111111111111111111000, 24'b111111111111110101001011, 24'b111111111111011110011110, 24'b000000000000011001100111, 24'b000000000000000000101100, 24'b000000000000100110100111, 24'b000000000000000000000000, 24'b111111111111111111111111, 24'b000000000000000110000101, 24'b111111111111100101001011, 24'b000000000000001110111110, 24'b000000000000000000000000, 24'b111111111111111001100010, 24'b111111111111101000110111, 24'b000000000000011000101111, 24'b111111111111111111111111, 24'b000000000000010110001101, 24'b000000000000001101110111, 24'b000000000000001101000011, 24'b111111111111111110110011, 24'b111111111111111111011110, 24'b111111111111001100010001, 24'b111111111111110111111011, 24'b111111111111111100010110, 24'b111111111111111111111110}, 
{24'b111111111111101101111001, 24'b111111111111101010100011, 24'b111111111111100100011000, 24'b111111111111111011100011, 24'b111111111111110111011110, 24'b000000000000000110101011, 24'b111111111111010011010100, 24'b111111111111110110011001, 24'b111111111111110001101001, 24'b111111111111111111111111, 24'b111111111111101101100110, 24'b000000000000010110010001, 24'b000000000000000010010001, 24'b000000000000001000110100, 24'b000000000000010011111101, 24'b000000000000000000000001, 24'b000000000000110011000001, 24'b000000000000000101101110, 24'b000000000000001111100010, 24'b000000000000010001001011, 24'b111111111111110101111110, 24'b000000000000010111010000, 24'b111111111111110000011110, 24'b111111111111011111111000, 24'b000000000000001011000110, 24'b000000000000100001000100, 24'b111111111111111111101110, 24'b000000000000000011011100, 24'b111111111111000011001001, 24'b000000000000010010010101, 24'b000000000000010001000110, 24'b111111111111101000000111, 24'b000000000000011110001011, 24'b000000000000101010100010, 24'b000000000000000000000000, 24'b000000000000010101111010, 24'b111111111111111111111111, 24'b000000000000010010001100, 24'b000000000000001100101111, 24'b000000000000000000000000, 24'b111111111111111000011101, 24'b111111111111101000101110, 24'b000000000000001001001011, 24'b000000000000011110111011, 24'b000000000000100001001110, 24'b111111111111110101001111, 24'b111111111111111010101010, 24'b111111111111110011110110, 24'b111111111111110111010110, 24'b000000000000000111100100, 24'b000000000000000000001101, 24'b000000000000000010001011, 24'b000000000000000000000000, 24'b000000000000001011100110, 24'b111111111111110100110101, 24'b000000000000110001010101, 24'b000000000000010110110010, 24'b111111111111111110011010, 24'b000000000000011000111110, 24'b000000000000001101111001, 24'b111111111110010111111111, 24'b111111111111011011000111, 24'b111111111111110100111110, 24'b111111111111111111010111}, 
{24'b000000000000000000010101, 24'b000000000000001111010011, 24'b111111111111111111111110, 24'b111111111111111111111101, 24'b111111111111101011011000, 24'b111111111111111110000000, 24'b111111111111101111100001, 24'b000000000000000000000000, 24'b000000000000000001110000, 24'b000000000000011000111000, 24'b000000000000000000111011, 24'b111111111111100111110100, 24'b111111111111111011111111, 24'b000000000000000000000000, 24'b111111111111111100101000, 24'b111111111111100011001110, 24'b111111111111001001101100, 24'b111111111111111111111110, 24'b111111111111011001010100, 24'b111111111111100011011101, 24'b111111111111100111000100, 24'b000000000000010110001110, 24'b000000000000000011000000, 24'b111111111111110110111000, 24'b111111111111100100000010, 24'b000000000000001001111100, 24'b000000000000000000000000, 24'b000000000000011111111101, 24'b000000000000110011100101, 24'b111111111111111101011011, 24'b000000000000000000000010, 24'b000000000000001110110000, 24'b111111111111010100010101, 24'b111111111111101000010000, 24'b000000000000000011100011, 24'b000000000000000101111011, 24'b111111111111101110000010, 24'b000000000000001111010101, 24'b000000000000001000011100, 24'b111111111111110110001110, 24'b111111111111100101001000, 24'b111111111111111101101000, 24'b000000000000000010000110, 24'b111111111111110101010111, 24'b000000000000000011100100, 24'b000000000000001110101011, 24'b111111111111111000010111, 24'b000000000000000001100001, 24'b000000000000000000000000, 24'b111111111111110010000011, 24'b111111111111100111001001, 24'b000000000000011010100111, 24'b000000000000001000000111, 24'b111111111111110100100110, 24'b000000000000001000011110, 24'b111111111111111100000011, 24'b111111111111100001101000, 24'b111111111111110111011110, 24'b111111111111111100101010, 24'b111111111111111011100000, 24'b000000000000110101001001, 24'b000000000000001100001101, 24'b111111111111111100111001, 24'b111111111111111111111110}, 
{24'b000000000000000000111100, 24'b000000000000100101100011, 24'b111111111111011010110101, 24'b111111111111110001001101, 24'b000000000000010100101001, 24'b111111111111110010110011, 24'b000000000001001101100001, 24'b111111111111101101100101, 24'b111111111111111111111111, 24'b000000000000010010110001, 24'b000000000000010000010001, 24'b111111111111111111110101, 24'b111111111111111100111011, 24'b111111111111100001001001, 24'b000000000000010010000000, 24'b000000000000001010001110, 24'b111111111111110011100110, 24'b111111111111111111111111, 24'b000000000000000000000000, 24'b000000000000000000000001, 24'b000000000000010000111110, 24'b111111111111100010100101, 24'b000000000000011001000110, 24'b000000000000100111001110, 24'b111111111111111010011010, 24'b111111111111111111111110, 24'b111111111111111110111101, 24'b111111111111111111111111, 24'b000000000000101111000111, 24'b000000000000000000010100, 24'b111111111111101110100000, 24'b000000000000000000000000, 24'b000000000000011000100101, 24'b111111111111001100000110, 24'b111111111111011101011001, 24'b000000000000001100101110, 24'b000000000000001000110111, 24'b111111111111011011011011, 24'b111111111111110011111001, 24'b111111111111110010010010, 24'b000000000000011001101010, 24'b000000000000011001000001, 24'b000000000000000000000000, 24'b111111111111101110101110, 24'b000000000000000000000011, 24'b000000000000011001010011, 24'b111111111111111100001110, 24'b111111111111111111111111, 24'b000000000000000000101111, 24'b000000000000001111101011, 24'b111111111111111100010100, 24'b111111111111110011100111, 24'b000000000000010110000001, 24'b111111111111110010001111, 24'b000000000000010001111001, 24'b000000000000100101011010, 24'b000000000000000010100011, 24'b000000000000010000110111, 24'b111111111111100110011000, 24'b111111111111101000100001, 24'b000000000000110101001111, 24'b111111111111110111110000, 24'b000000000000000010111100, 24'b111111111111111010000001}, 
{24'b000000000000000001000010, 24'b111111111111100011000010, 24'b000000000000010111100110, 24'b111111111111101101110101, 24'b111111111111111111110011, 24'b000000000000001101100010, 24'b111111111111011010110000, 24'b000000000000001100010000, 24'b000000000000011111011001, 24'b000000000000001001110111, 24'b000000000000010111001100, 24'b000000000000010100101001, 24'b111111111111101100011111, 24'b111111111111111011001001, 24'b111111111111111100101101, 24'b000000000000000000000100, 24'b111111111111000010100101, 24'b000000000000010100101011, 24'b111111111111111101101011, 24'b000000000000000001111111, 24'b111111111111101001011100, 24'b000000000000000100011110, 24'b000000000000001001110011, 24'b111111111111111111111110, 24'b111111111111100010100010, 24'b111111111111111100111100, 24'b111111111111111010110000, 24'b000000000001001111110111, 24'b111111111111010101100110, 24'b000000000000000100010000, 24'b000000000000000110001101, 24'b111111111111111100010000, 24'b111111111111110001110111, 24'b000000000000000111011101, 24'b111111111111111010111111, 24'b111111111111110111011001, 24'b111111111111110100100110, 24'b111111111111110010100011, 24'b111111111111111110100101, 24'b111111111111101100111101, 24'b000000000000010100100110, 24'b000000000000000111111001, 24'b000000000000011111110010, 24'b000000000000000101100111, 24'b000000000000000010010111, 24'b111111111111101101011000, 24'b000000000000000000000000, 24'b111111111111111111111111, 24'b111111111111111111111110, 24'b000000000000001100011001, 24'b000000000000001011010110, 24'b000000000000010010110111, 24'b111111111111111111100111, 24'b111111111111101101001110, 24'b000000000000000000100100, 24'b000000000000000000000000, 24'b000000000000010100101000, 24'b111111111111110011001001, 24'b111111111111011100110001, 24'b000000000000100011111011, 24'b111111111111101101001100, 24'b000000000001001010011111, 24'b111111111111111110101110, 24'b111111111111101001010100}, 
{24'b111111111111011011000111, 24'b111111111111111111111000, 24'b111111111111100101110010, 24'b000000000000001110101111, 24'b000000000000010000110110, 24'b111111111111111001011100, 24'b000000000000100001000101, 24'b111111111111110101000110, 24'b111111111111100001010100, 24'b111111111111101000100001, 24'b111111111111101111111011, 24'b111111111111100001100010, 24'b111111111111110001010110, 24'b000000000000001100100110, 24'b000000000000000000000000, 24'b000000000000000000000001, 24'b000000000000110101111011, 24'b111111111111111101001111, 24'b111111111111111111111011, 24'b000000000000011010010100, 24'b000000000000010010101111, 24'b111111111111011010111101, 24'b111111111111100111100001, 24'b000000000000001100000110, 24'b111111111111100100011100, 24'b111111111111111110101010, 24'b111111111111101111011000, 24'b111111111111101010100111, 24'b111111111111100100000111, 24'b000000000000010011010101, 24'b000000000000001110100101, 24'b111111111111110110000001, 24'b111111111111111011010110, 24'b111111111111000001101010, 24'b111111111111110100101100, 24'b000000000000000011001010, 24'b111111111111110111101101, 24'b111111111111101101000001, 24'b111111111111111111110001, 24'b000000000000000111100111, 24'b111111111111111000011000, 24'b111111111111111111110101, 24'b111111111111111101110000, 24'b111111111111010101011111, 24'b000000000000000000000011, 24'b000000000000000000000000, 24'b000000000000010101110001, 24'b111111111111111000000010, 24'b000000000000011011000111, 24'b111111111111110011110011, 24'b000000000000010010011011, 24'b111111111111111111111010, 24'b000000000000001110011100, 24'b111111111111100110111101, 24'b111111111111111111111111, 24'b000000000000100000110001, 24'b000000000000010100000000, 24'b000000000000010010101100, 24'b000000000000000001100111, 24'b111111111111100110011010, 24'b111111111111101100110111, 24'b111111111111010100000101, 24'b111111111111111111111000, 24'b000000000000000110110110}, 
{24'b000000000000010011101111, 24'b000000000000000000001010, 24'b000000000000001000011001, 24'b111111111111111111111111, 24'b000000000000001001110100, 24'b111111111111110111011000, 24'b000000000000001111000001, 24'b000000000000000010101101, 24'b000000000000001000101100, 24'b000000000000010101110000, 24'b111111111111101111001000, 24'b111111111111111110101011, 24'b111111111111111111011110, 24'b111111111111111111011100, 24'b111111111111010101110001, 24'b111111111111101100111100, 24'b000000000000101000010110, 24'b111111111111111110001101, 24'b111111111111111100101010, 24'b000000000000000000000001, 24'b111111111111100111101010, 24'b000000000000000000100101, 24'b000000000000010000000011, 24'b000000000000000010011011, 24'b000000000000000010010110, 24'b000000000000010101101010, 24'b000000000000000000000000, 24'b000000000000000010011010, 24'b000000000000000000000000, 24'b111111111111111100111110, 24'b111111111111110011001001, 24'b111111111111010101011000, 24'b000000000000010000111010, 24'b000000000000010101111100, 24'b111111111111111110001000, 24'b111111111111110000111110, 24'b000000000000000000000000, 24'b111111111111010110000110, 24'b111111111111111101000100, 24'b111111111111111111110010, 24'b000000000000001100100010, 24'b111111111111110111101001, 24'b111111111111111111111111, 24'b000000000000110110001110, 24'b000000000000011100101100, 24'b111111111111111111100111, 24'b111111111111111111111110, 24'b111111111111111111111111, 24'b111111111111110000100110, 24'b000000000000001001011010, 24'b000000000000001001001110, 24'b000000000000001011001011, 24'b000000000000001010000100, 24'b000000000000011000110110, 24'b000000000000010110011000, 24'b000000000000101010001101, 24'b111111111111110111000011, 24'b000000000000011001001011, 24'b000000000000001001110001, 24'b111111111111101011001001, 24'b000000000000000111000110, 24'b111111111111100111001001, 24'b111111111111100011110110, 24'b111111111111100000000101}, 
{24'b000000000000000000000001, 24'b000000000000001110100111, 24'b111111111111110011100010, 24'b000000000000000000000000, 24'b111111111111111100110111, 24'b111111111111111101110100, 24'b111111111111010101101110, 24'b111111111111111111111111, 24'b000000000000010000001110, 24'b000000000000001111111111, 24'b000000000000001111001101, 24'b111111111111100110100001, 24'b111111111111111010010010, 24'b000000000000010010001011, 24'b111111111111111111111110, 24'b000000000000000000010011, 24'b111111111111001010001001, 24'b111111111111111111111110, 24'b000000000000010111110101, 24'b000000000000000100100000, 24'b000000000000001111001111, 24'b111111111111111000100111, 24'b000000000000001111111110, 24'b000000000000011001111010, 24'b111111111111101001010000, 24'b111111111111101110000110, 24'b111111111111111111101011, 24'b111111111111111010110101, 24'b000000000000000100010011, 24'b000000000000000000000000, 24'b111111111111111111111111, 24'b000000000000010100000111, 24'b111111111111010000000000, 24'b000000000000010111001000, 24'b000000000000100000000101, 24'b000000000000000111011101, 24'b000000000000000111001100, 24'b111111111111111001000101, 24'b000000000000000111010111, 24'b111111111111111001001010, 24'b111111111111101111111011, 24'b111111111111111100110001, 24'b000000000000001010100001, 24'b000000000000101100110000, 24'b111111111111001001110000, 24'b111111111111100011011110, 24'b000000000000001100010010, 24'b111111111111111001101111, 24'b000000000000011100110101, 24'b111111111111110000111000, 24'b111111111111101010110100, 24'b111111111111101110000100, 24'b111111111111111111111111, 24'b000000000000000111101100, 24'b111111111111110101111011, 24'b111111111111001010011101, 24'b111111111111110110110110, 24'b111111111111111111010110, 24'b000000000000000010110010, 24'b111111111111011000111100, 24'b000000000001000111101011, 24'b111111111111011101001010, 24'b000000000000100010101010, 24'b000000000000001001110011}, 
{24'b000000000000000101000000, 24'b111111111111110011101110, 24'b000000000000101000001101, 24'b111111111111101100101001, 24'b111111111111100010010110, 24'b000000000000000101110000, 24'b000000000000010011110011, 24'b000000000000010011001111, 24'b111111111111110100101001, 24'b111111111111110101101110, 24'b000000000000000011010111, 24'b000000000000001110101010, 24'b000000000000001111000010, 24'b000000000000000011001101, 24'b111111111111110010111011, 24'b000000000000001000001110, 24'b000000000000011110001000, 24'b111111111111111111010010, 24'b111111111111101110000110, 24'b000000000000000000000000, 24'b000000000000000100110000, 24'b000000000000000001010011, 24'b111111111111101101001111, 24'b000000000000000111001110, 24'b000000000000110010010111, 24'b000000000000000000101001, 24'b000000000000001011100011, 24'b111111111111001101001111, 24'b111111111111111011010110, 24'b000000000000000000100110, 24'b111111111111110011011100, 24'b111111111111101100000011, 24'b000000000000011101010101, 24'b111111111111111110010011, 24'b111111111111111101100101, 24'b111111111111101100011110, 24'b000000000000001000110111, 24'b000000000000010010101100, 24'b111111111111111111011000, 24'b111111111111111101001110, 24'b111111111111110100000011, 24'b000000000000001110100111, 24'b000000000000000000000000, 24'b111111111111010100000100, 24'b000000000000010011111010, 24'b000000000000011001100010, 24'b111111111111111111111111, 24'b000000000000000001101000, 24'b111111111111100100001110, 24'b111111111111111011001101, 24'b111111111111111111111111, 24'b111111111111101011101011, 24'b000000000000000000000000, 24'b111111111111110100111100, 24'b000000000000000011101010, 24'b111111111111001011101100, 24'b111111111111111111111111, 24'b111111111111111111111100, 24'b000000000000010001100111, 24'b000000000000100100000010, 24'b111111111111010011100001, 24'b000000000000100001010010, 24'b000000000000000010010111, 24'b111111111111111011001110}, 
{24'b000000000000010010011010, 24'b000000000001001111011000, 24'b000000000000011111101101, 24'b000000000000010010010000, 24'b111111111111100001011011, 24'b111111111111101011101011, 24'b111111111101011001101000, 24'b111111111111100010110000, 24'b000000000000011001110010, 24'b111111111111111111111111, 24'b000000000000010010110100, 24'b000000000000110111001111, 24'b000000000000000100011100, 24'b000000000000000000010110, 24'b111111111111111110111010, 24'b000000000000000000000000, 24'b111111111111110011111000, 24'b111111111111110011000010, 24'b000000000000001110101110, 24'b111111111111011111110111, 24'b111111111111010101011100, 24'b111111111111111001011011, 24'b111111111111011010101000, 24'b000000000000000001111000, 24'b111111111101101110010011, 24'b000000000000110100001011, 24'b000000000000111111010011, 24'b000000000000100110101000, 24'b111111111110010000011011, 24'b111111111111101011111110, 24'b111111111111010011111110, 24'b111111111111001010000000, 24'b111111111101011110011001, 24'b000000000000101011010010, 24'b111111111111111101001100, 24'b000000000000010100011001, 24'b000000000000000001100001, 24'b111111111110100100010010, 24'b000000000000000000000001, 24'b000000000000000000000000, 24'b000000000000000010000010, 24'b000000000001000001001111, 24'b111111111111110010111000, 24'b111111111111010110101110, 24'b000000000000111001011011, 24'b111111111111100011100110, 24'b111111111111101011001111, 24'b111111111111100110111000, 24'b000000000000011110100011, 24'b000000000000100010000000, 24'b111111111111111011101001, 24'b111111111111101001101010, 24'b111111111111111111110111, 24'b111111111111111000110011, 24'b000000000000000000000000, 24'b111111111111100111110111, 24'b000000000000100110110100, 24'b000000000001000101011001, 24'b000000000000101101100010, 24'b111111111111000101110101, 24'b111111111100010011000000, 24'b000000000000111000101010, 24'b000000000000000101111010, 24'b000000000000010100010010}, 
{24'b111111111111110000100010, 24'b000000000000010101100101, 24'b000000000000010100010100, 24'b111111111111111111111001, 24'b111111111111101000001100, 24'b111111111111111010010000, 24'b111111111111100111011100, 24'b111111111111111100011100, 24'b000000000000001001100010, 24'b111111111111111011001100, 24'b111111111111111110000001, 24'b111111111111111101011111, 24'b111111111111111111111101, 24'b111111111111110100010001, 24'b111111111111111110010010, 24'b111111111111111001100101, 24'b000000000000010100000011, 24'b111111111111111111111111, 24'b111111111111010110111110, 24'b000000000000011101110000, 24'b000000000000100110000110, 24'b000000000000011010100010, 24'b111111111111101011101101, 24'b111111111111110111001110, 24'b111111111111101001110111, 24'b111111111111101101011100, 24'b000000000000001110100001, 24'b000000000000001110111110, 24'b000000000000001110011110, 24'b000000000000010111000001, 24'b000000000000000010001100, 24'b000000000000011000101101, 24'b111111111111111101010100, 24'b000000000000000000010011, 24'b000000000000010011011111, 24'b000000000000001000011010, 24'b111111111111111011110001, 24'b111111111111111111011001, 24'b000000000000000000000000, 24'b111111111111101101010001, 24'b111111111111110001101101, 24'b111111111111111000111100, 24'b111111111111101001000001, 24'b000000000000011100110010, 24'b000000000000000000000001, 24'b111111111111111111101001, 24'b111111111111111010101101, 24'b111111111111110110100011, 24'b111111111111001100011100, 24'b111111111111111101100001, 24'b111111111111110001101000, 24'b111111111111110110111011, 24'b111111111111111001100110, 24'b000000000000010000111011, 24'b000000000000101011101001, 24'b000000000000001011111111, 24'b111111111111111111001001, 24'b111111111111101010000011, 24'b111111111111111110000111, 24'b000000000000000000000001, 24'b000000000000010100110101, 24'b111111111111111110101001, 24'b000000000000000010111011, 24'b000000000000000000000000}
};

localparam logic signed [23:0] bias [64] = '{
24'b111111111111111101100111,  // -0.037350185215473175
24'b000000000000010001100000,  // 0.27355897426605225
24'b111111111111111000000100,  // -0.12378914654254913
24'b111111111111111011110111,  // -0.064457006752491
24'b000000000000000011011111,  // 0.05452875792980194
24'b000000000000000111011110,  // 0.11671770364046097
24'b000000000000001000101110,  // 0.13640816509723663
24'b000000000000000100110010,  // 0.07482525706291199
24'b000000000000000010111111,  // 0.04674031585454941
24'b111111111111110011000110,  // -0.20146161317825317
24'b111111111111111001101010,  // -0.09910125285387039
24'b000000000000001001101010,  // 0.15104414522647858
24'b111111111111111001011101,  // -0.10221704095602036
24'b111111111111110110101001,  // -0.1461549550294876
24'b111111111111111010011110,  // -0.08641516417264938
24'b000000000000001010101000,  // 0.16613510251045227
24'b111111111111111010101001,  // -0.0836295336484909
24'b111111111111111100010100,  // -0.05756539851427078
24'b111111111111111101111011,  // -0.03229188174009323
24'b111111111111111110001011,  // -0.028388574719429016
24'b000000000000001000000100,  // 0.1260243058204651
24'b111111111111111101101000,  // -0.037064336240291595
24'b000000000000001100011000,  // 0.19336333870887756
24'b000000000000000001010111,  // 0.02124214917421341
24'b000000000000011111111010,  // 0.4985624849796295
24'b000000000000000001000000,  // 0.0158411655575037
24'b111111111111111010101100,  // -0.08296407759189606
24'b000000000000000111000100,  // 0.11056788265705109
24'b000000000000000000110000,  // 0.01173810102045536
24'b111111111111111001000011,  // -0.10843746364116669
24'b000000000000010001100011,  // 0.27439257502555847
24'b000000000000000101111000,  // 0.09199801832437515
24'b000000000000010001100011,  // 0.27419957518577576
24'b000000000000010001010100,  // 0.27063727378845215
24'b111111111111110000000111,  // -0.24828937649726868
24'b000000000000000101000000,  // 0.07818280160427094
24'b111111111111111111101000,  // -0.005749030504375696
24'b000000000000000110111100,  // 0.10850494354963303
24'b000000000000001000101100,  // 0.13591453433036804
24'b111111111111111000010000,  // -0.12088628858327866
24'b111111111111111100010111,  // -0.05666546896100044
24'b000000000000000101111101,  // 0.09311636537313461
24'b000000000000000011100000,  // 0.05477767437696457
24'b000000000000000001111001,  // 0.029585206881165504
24'b111111111111101100000001,  // -0.31209176778793335
24'b111111111111111010100101,  // -0.08465463668107986
24'b111111111111110101010000,  // -0.16775836050510406
24'b000000000000001001011100,  // 0.14762157201766968
24'b111111111111110000111000,  // -0.23618532717227936
24'b000000000000000100001011,  // 0.06535740196704865
24'b111111111111110111110001,  // -0.12853026390075684
24'b111111111111110111001010,  // -0.13802281022071838
24'b111111111111110110010011,  // -0.15156887471675873
24'b000000000000000101000110,  // 0.07979883998632431
24'b000000000000001011100111,  // 0.18141601979732513
24'b111111111111111100100010,  // -0.054039113223552704
24'b111111111111111111010110,  // -0.010052933357656002
24'b000000000000000100001110,  // 0.06611225008964539
24'b000000000000000011001110,  // 0.05053366720676422
24'b000000000000000001101110,  // 0.026860840618610382
24'b000000000000000010000110,  // 0.03283466026186943
24'b000000000000001001111101,  // 0.15558314323425293
24'b111111111111101101101011,  // -0.2863388657569885
24'b111111111111111010011000   // -0.08769102394580841
};
endpackage