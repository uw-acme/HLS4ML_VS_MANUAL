// Width: 16
// NFRAC: 10
package dense_4_16_10;

localparam logic signed [15:0] weights [32][5] = '{ 
{16'b1111111111110011, 16'b0000000101000011, 16'b1111111011001110, 16'b0000000001000011, 16'b1111111110010011}, 
{16'b1111110111000100, 16'b1111111111000111, 16'b0000000111010111, 16'b1111111111110011, 16'b0000000000010001}, 
{16'b0000000101111100, 16'b0000000011011000, 16'b1111111111100011, 16'b1111111001100000, 16'b1111111100101000}, 
{16'b1111111001111111, 16'b1111111010000010, 16'b1111111110001101, 16'b0000000100111011, 16'b0000000011110000}, 
{16'b0000000001111101, 16'b0000000010000011, 16'b0000000010100000, 16'b1111111111101101, 16'b1111101111110010}, 
{16'b0000000101001110, 16'b1111111001101100, 16'b0000000010111001, 16'b1111111101011010, 16'b1111111101010001}, 
{16'b1111111001100101, 16'b0000000000100100, 16'b1111111111111111, 16'b0000000010110010, 16'b0000000001000110}, 
{16'b1111111111111110, 16'b0000000100100011, 16'b1111111001101110, 16'b0000000010100110, 16'b0000000010001011}, 
{16'b0000000010100111, 16'b1111111101010010, 16'b0000000000000001, 16'b1111111000100111, 16'b1111111100000001}, 
{16'b1111111111111111, 16'b1111111011101111, 16'b0000000010110110, 16'b0000000110111000, 16'b0000000000000000}, 
{16'b1111111101111010, 16'b1111111101101011, 16'b0000000000000000, 16'b0000001001010011, 16'b1111111011101101}, 
{16'b0000000010101101, 16'b0000000011101010, 16'b1111111010100011, 16'b1111111111100011, 16'b0000000001111100}, 
{16'b0000000000000000, 16'b0000000010101011, 16'b0000000000001001, 16'b1111111100101011, 16'b1111110110000010}, 
{16'b0000000010110101, 16'b0000000001000001, 16'b0000000110101101, 16'b1111111110111000, 16'b1111111001001001}, 
{16'b0000000001011100, 16'b1111111111001110, 16'b1111111010001110, 16'b1111111111011110, 16'b0000001000100101}, 
{16'b1111111000011010, 16'b1111111100000101, 16'b1111111100011100, 16'b0000000110011000, 16'b0000000000100000}, 
{16'b0000000101100010, 16'b1111111101010000, 16'b1111111101110101, 16'b1111111100011000, 16'b1111111111000010}, 
{16'b0000000011000111, 16'b1111111111010110, 16'b1111111001011001, 16'b1111111111100000, 16'b0000000001001000}, 
{16'b0000000100001000, 16'b0000000000101010, 16'b1111111100100000, 16'b0000000000000000, 16'b1111111001111111}, 
{16'b0000000011101100, 16'b1111111110100111, 16'b1111111100100110, 16'b0000000011010100, 16'b0000000001100001}, 
{16'b0000000001000101, 16'b1111111111100000, 16'b0000000100110000, 16'b1111111001000110, 16'b1111111111101010}, 
{16'b0000000000000000, 16'b0000000001111000, 16'b0000000111110010, 16'b1111110111101101, 16'b1111110110000111}, 
{16'b1111111110011011, 16'b0000000001110000, 16'b0000000010110101, 16'b1111111010010010, 16'b0000001000010110}, 
{16'b1111111111111111, 16'b0000000010101000, 16'b0000000100100001, 16'b0000000000100110, 16'b1111110110110110}, 
{16'b1111111101010010, 16'b0000000101110101, 16'b1111111100011011, 16'b0000000000000101, 16'b0000000110001101}, 
{16'b0000000000011010, 16'b0000000100010000, 16'b0000000000011110, 16'b1111110100000010, 16'b0000001000110001}, 
{16'b1111111000101001, 16'b1111111100000110, 16'b0000000011011011, 16'b0000000011111010, 16'b0000000011001110}, 
{16'b0000000000000100, 16'b0000000011110110, 16'b1111111111011010, 16'b1111111101100101, 16'b0000000000100000}, 
{16'b1111111110010101, 16'b0000000011111100, 16'b1111110111111100, 16'b0000000010001110, 16'b1111111101011101}, 
{16'b1111111111101101, 16'b0000000010010000, 16'b1111111101010011, 16'b1111111001100101, 16'b0000001001011111}, 
{16'b0000000111001011, 16'b0000000001000111, 16'b0000000101001100, 16'b1111110110100100, 16'b1111111010111101}, 
{16'b1111111111000011, 16'b1111111001110100, 16'b0000000101110110, 16'b0000000001001000, 16'b0000000010000010}
};

localparam logic signed [15:0] bias [5] = '{
16'b1111111111000000,  // -0.06223141402006149
16'b1111111110111111,  // -0.06270556896924973
16'b1111111110111000,  // -0.07014333456754684
16'b0000000001010100,  // 0.0820775106549263
16'b0000000011011100   // 0.2155742198228836
};
endpackage