// Width: 14
// NFRAC: 7
package dense_4_14_7;

localparam logic signed [13:0] weights [32][5] = '{ 
{14'b11111111111110, 14'b00000000101000, 14'b11111111011001, 14'b00000000001000, 14'b11111111110010}, 
{14'b11111110111000, 14'b11111111111000, 14'b00000000111010, 14'b11111111111110, 14'b00000000000010}, 
{14'b00000000101111, 14'b00000000011011, 14'b11111111111100, 14'b11111111001100, 14'b11111111100101}, 
{14'b11111111001111, 14'b11111111010000, 14'b11111111110001, 14'b00000000100111, 14'b00000000011110}, 
{14'b00000000001111, 14'b00000000010000, 14'b00000000010100, 14'b11111111111101, 14'b11111101111110}, 
{14'b00000000101001, 14'b11111111001101, 14'b00000000010111, 14'b11111111101011, 14'b11111111101010}, 
{14'b11111111001100, 14'b00000000000100, 14'b11111111111111, 14'b00000000010110, 14'b00000000001000}, 
{14'b11111111111111, 14'b00000000100100, 14'b11111111001101, 14'b00000000010100, 14'b00000000010001}, 
{14'b00000000010100, 14'b11111111101010, 14'b00000000000000, 14'b11111111000100, 14'b11111111100000}, 
{14'b11111111111111, 14'b11111111011101, 14'b00000000010110, 14'b00000000110111, 14'b00000000000000}, 
{14'b11111111101111, 14'b11111111101101, 14'b00000000000000, 14'b00000001001010, 14'b11111111011101}, 
{14'b00000000010101, 14'b00000000011101, 14'b11111111010100, 14'b11111111111100, 14'b00000000001111}, 
{14'b00000000000000, 14'b00000000010101, 14'b00000000000001, 14'b11111111100101, 14'b11111110110000}, 
{14'b00000000010110, 14'b00000000001000, 14'b00000000110101, 14'b11111111110111, 14'b11111111001001}, 
{14'b00000000001011, 14'b11111111111001, 14'b11111111010001, 14'b11111111111011, 14'b00000001000100}, 
{14'b11111111000011, 14'b11111111100000, 14'b11111111100011, 14'b00000000110011, 14'b00000000000100}, 
{14'b00000000101100, 14'b11111111101010, 14'b11111111101110, 14'b11111111100011, 14'b11111111111000}, 
{14'b00000000011000, 14'b11111111111010, 14'b11111111001011, 14'b11111111111100, 14'b00000000001001}, 
{14'b00000000100001, 14'b00000000000101, 14'b11111111100100, 14'b00000000000000, 14'b11111111001111}, 
{14'b00000000011101, 14'b11111111110100, 14'b11111111100100, 14'b00000000011010, 14'b00000000001100}, 
{14'b00000000001000, 14'b11111111111100, 14'b00000000100110, 14'b11111111001000, 14'b11111111111101}, 
{14'b00000000000000, 14'b00000000001111, 14'b00000000111110, 14'b11111110111101, 14'b11111110110000}, 
{14'b11111111110011, 14'b00000000001110, 14'b00000000010110, 14'b11111111010010, 14'b00000001000010}, 
{14'b11111111111111, 14'b00000000010101, 14'b00000000100100, 14'b00000000000100, 14'b11111110110110}, 
{14'b11111111101010, 14'b00000000101110, 14'b11111111100011, 14'b00000000000000, 14'b00000000110001}, 
{14'b00000000000011, 14'b00000000100010, 14'b00000000000011, 14'b11111110100000, 14'b00000001000110}, 
{14'b11111111000101, 14'b11111111100000, 14'b00000000011011, 14'b00000000011111, 14'b00000000011001}, 
{14'b00000000000000, 14'b00000000011110, 14'b11111111111011, 14'b11111111101100, 14'b00000000000100}, 
{14'b11111111110010, 14'b00000000011111, 14'b11111110111111, 14'b00000000010001, 14'b11111111101011}, 
{14'b11111111111101, 14'b00000000010010, 14'b11111111101010, 14'b11111111001100, 14'b00000001001011}, 
{14'b00000000111001, 14'b00000000001000, 14'b00000000101001, 14'b11111110110100, 14'b11111111010111}, 
{14'b11111111111000, 14'b11111111001110, 14'b00000000101110, 14'b00000000001001, 14'b00000000010000}
};

localparam logic signed [13:0] bias [5] = '{
14'b11111111111000,  // -0.06223141402006149
14'b11111111110111,  // -0.06270556896924973
14'b11111111110111,  // -0.07014333456754684
14'b00000000001010,  // 0.0820775106549263
14'b00000000011011   // 0.2155742198228836
};
endpackage