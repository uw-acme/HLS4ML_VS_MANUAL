// Width: 27
// NFRAC: 13
package dense_2_27_14;

localparam logic signed [26:0] weights [64][32] = '{ 
{27'b000000000000000100010011011, 27'b000000000000000000001000010, 27'b111111111111111100111101100, 27'b111111111111111111101010011, 27'b000000000000000100001011011, 27'b000000000000000000000000000, 27'b111111111111111101101100001, 27'b111111111111111111111111111, 27'b111111111111111011100111100, 27'b000000000000000001010001101, 27'b000000000000000000000000000, 27'b111111111111111111111010001, 27'b111111111111111111111111100, 27'b111111111111111100110011001, 27'b111111111111111111001100001, 27'b111111111111111011110011111, 27'b000000000000000000000000000, 27'b111111111111111111110010101, 27'b111111111111111100111100111, 27'b111111111111111101011101110, 27'b000000000000000000000000000, 27'b000000000000000000000000000, 27'b111111111111111111110111110, 27'b111111111111111111111101001, 27'b000000000000000000000000000, 27'b000000000000000001100110111, 27'b000000000000000110001011010, 27'b000000000000000010110011011, 27'b111111111111111111111111100, 27'b000000000000000000110011110, 27'b111111111111111001011100110, 27'b000000000000000000000000010}, 
{27'b111111111111111110011001011, 27'b111111111111111101100001011, 27'b111111111111111101110010010, 27'b111111111111111111000111001, 27'b111111111111111111111010001, 27'b000000000000000000101100000, 27'b111111111111111100011011010, 27'b000000000000000000000101011, 27'b000000000000000000000100111, 27'b111111111111111110111111100, 27'b000000000000000010011111111, 27'b111111111111111111010011100, 27'b111111111111111111000011101, 27'b111111111111111100100001111, 27'b000000000000000000000111101, 27'b111111111111111111001110110, 27'b000000000000000000001100110, 27'b111111111111111100111000100, 27'b000000000000000010101111111, 27'b000000000000000011101011000, 27'b111111111111111111011111111, 27'b111111111111111111111010001, 27'b111111111111111111111111101, 27'b000000000000000000011000001, 27'b111111111111111110110111000, 27'b000000000000000100011001101, 27'b000000000000000011111101100, 27'b000000000000000000001000101, 27'b000000000000000000011101001, 27'b111111111111111000001101100, 27'b000000000000000000000111100, 27'b000000000000000000000000000}, 
{27'b000000000000000001001010001, 27'b111111111111111110001010100, 27'b111111111111111101111011010, 27'b111111111111111111010101001, 27'b111111111111111110110000101, 27'b111111111111111110101000101, 27'b111111111111111101000010101, 27'b000000000000000000000100100, 27'b111111111111111101110101110, 27'b000000000000000000001001001, 27'b000000000000000000000010001, 27'b111111111111111110101101011, 27'b000000000000000001011100100, 27'b111111111111111110111101111, 27'b111111111111111111111110100, 27'b111111111111111111011010011, 27'b000000000000000000000101000, 27'b000000000000000001100001110, 27'b000000000000000000111100000, 27'b000000000000000011101011010, 27'b000000000000000000101010000, 27'b111111111111111110101001111, 27'b000000000000000000000000011, 27'b000000000000000000100011110, 27'b111111111111111111101101001, 27'b000000000000000011010110010, 27'b000000000000000010011000110, 27'b000000000000000001100011001, 27'b111111111111111111111111100, 27'b111111111111111101100100010, 27'b111111111111111111110010001, 27'b000000000000000001100101101}, 
{27'b000000000000000010001101011, 27'b000000000000000000010011101, 27'b000000000000000000110110001, 27'b111111111111111111110110000, 27'b111111111111110111110110101, 27'b000000000000000000000000000, 27'b000000000000000000000000010, 27'b000000000000000011100111100, 27'b000000000000000011111000011, 27'b111111111111111111110010011, 27'b111111111111111111111111111, 27'b000000000000000000000000000, 27'b000000000000000000000000010, 27'b000000000000000000000101000, 27'b111111111111111111101101010, 27'b000000000000000011011011111, 27'b000000000000000000000000001, 27'b111111111111111111100110110, 27'b111111111111111111111111111, 27'b111111111111111101001011101, 27'b111111111111111111000001010, 27'b000000000000000000110010101, 27'b111111111111111110111111000, 27'b111111111111111111111111101, 27'b000000000000000000000011111, 27'b111111111111111111001100000, 27'b000000000000000001001010110, 27'b111111111111111111111111110, 27'b111111111111111111111111111, 27'b111111111111111111111111111, 27'b111111111111111100100011101, 27'b000000000000000100111101101}, 
{27'b111111111111110101000101001, 27'b111111111111111111100110100, 27'b111111111111111111111011101, 27'b000000000000000000000101011, 27'b111111111111111111100101000, 27'b000000000000000000000110110, 27'b111111111111111111001101101, 27'b111111111111111101100110101, 27'b000000000000000000110111100, 27'b111111111111111111101011010, 27'b111111111111111111110010000, 27'b111111111111111111111111110, 27'b111111111111111111111111110, 27'b000000000000000011010111010, 27'b000000000000000000000000000, 27'b000000000000000101010000111, 27'b111111111111111111111111111, 27'b000000000000000011011111011, 27'b111111111111111001100110011, 27'b000000000000000000000000010, 27'b111111111111111110001101101, 27'b000000000000000010101100100, 27'b000000000000000100001000011, 27'b000000000000000000000000000, 27'b000000000000000000101110011, 27'b000000000000000010100110110, 27'b000000000000000011110100011, 27'b000000000000000000010001110, 27'b111111111111111111111011011, 27'b111111111111111111111111110, 27'b111111111111111111110001111, 27'b000000000000000011100111101}, 
{27'b000000000000000000111011000, 27'b111111111111111111111111110, 27'b000000000000000010011000110, 27'b111111111111110101100111111, 27'b111111111111101001111101110, 27'b111111111111111010011001001, 27'b000000000000000101101010101, 27'b111111111111110110000010111, 27'b111111111111111111111111101, 27'b111111111111110101001010011, 27'b111111111111110111111110111, 27'b111111111111111010100010110, 27'b000000000000000101101001110, 27'b111111111111111111111111111, 27'b111111111111111111110000110, 27'b000000000000000000000000000, 27'b111111111111111111111111111, 27'b111111111111111111111111100, 27'b111111111111111101111000100, 27'b111111111111111111111111111, 27'b111111111111111000001011000, 27'b000000000000000000000000000, 27'b000000000000000010111110011, 27'b111111111111111111111111111, 27'b000000000000000000010110100, 27'b000000000000000100010010001, 27'b000000000000000000110100011, 27'b111111111111111111111111111, 27'b111111111111111111111111111, 27'b000000000000000011010010100, 27'b111111111111111111011101000, 27'b000000000000000011001101011}, 
{27'b111111111111111111011011001, 27'b111111111111111101011110111, 27'b111111111111111100001000100, 27'b111111111111111111001111111, 27'b111111111111111011011000100, 27'b000000000000000001000011101, 27'b111111111111111101000111101, 27'b111111111111111101101110100, 27'b111111111111111001010111010, 27'b000000000000000000110001100, 27'b111111111111111111111010110, 27'b111111111111111101011101000, 27'b000000000000000001111001110, 27'b111111111111111111110101101, 27'b111111111111111111010101100, 27'b111111111111110111001001000, 27'b111111111111111111111111110, 27'b000000000000000001010110000, 27'b000000000000000011000100010, 27'b111111111111111101011001110, 27'b111111111111111101100110011, 27'b111111111111111110111111111, 27'b111111111111111111111110101, 27'b000000000000000000011100010, 27'b111111111111111111010001011, 27'b111111111111110101101000010, 27'b111111111111111011110000101, 27'b111111111111111111010001111, 27'b000000000000000000000101110, 27'b111111111111111111101010001, 27'b000000000000000000011111010, 27'b111111111111111111111111010}, 
{27'b111111111111111101100010110, 27'b111111111111111110100011011, 27'b111111111111111110101110101, 27'b111111111111111100001101000, 27'b111111111111111110001001011, 27'b111111111111111111111111101, 27'b000000000000000001101010111, 27'b111111111111111110101111000, 27'b000000000000000011001101011, 27'b000000000000000000000000001, 27'b000000000000000000000000000, 27'b111111111111111111111111111, 27'b000000000000000011100000000, 27'b000000000000000000000000001, 27'b111111111111111111111111110, 27'b111111111111111110110111100, 27'b111111111111111111111111100, 27'b000000000000000000000000000, 27'b111111111111111111111111100, 27'b000000000000000000000000000, 27'b111111111111111111111111101, 27'b111111111111111111111111011, 27'b000000000000000000000000001, 27'b111111111111111111111111111, 27'b000000000000000000101101001, 27'b111111111111111101000111101, 27'b000000000000000000001110001, 27'b111111111111111111111111101, 27'b111111111111111110110110001, 27'b111111111111111111111111010, 27'b000000000000000000000000011, 27'b111111111111111111111111110}, 
{27'b111111111111111000010111000, 27'b111111111111111111000101100, 27'b111111111111111001111010110, 27'b000000000000000001111101001, 27'b000000000000000111110010101, 27'b111111111111111111111111111, 27'b111111111111111111100010010, 27'b000000000000000011110100101, 27'b111111111111111000111110101, 27'b111111111111111111010000001, 27'b000000000000000000000000000, 27'b111111111111111100110001101, 27'b111111111111111111111111101, 27'b000000000000000001001101111, 27'b111111111111111100111100111, 27'b000000000000001100000100000, 27'b111111111111111111110111001, 27'b000000000000000000101111111, 27'b000000000000000011010100101, 27'b000000000000000011111010110, 27'b000000000000000000000000001, 27'b111111111111111010101000001, 27'b000000000000000000000000001, 27'b000000000000000110100101011, 27'b111111111111111101000110011, 27'b000000000000001011001010011, 27'b111111111111111101100111001, 27'b111111111111111100101111001, 27'b111111111111111000011100101, 27'b111111111111111000100100101, 27'b000000000000000000000000010, 27'b000000000000000000110110101}, 
{27'b000000000000000000000000001, 27'b111111111111111111110000001, 27'b111111111111111110110100011, 27'b000000000000000000000000000, 27'b000000000000000100111011111, 27'b111111111111111111101011010, 27'b111111111111111110111110110, 27'b000000000000000001011110000, 27'b000000000000000001100111111, 27'b000000000000000000000011100, 27'b111111111111111111110111010, 27'b111111111111111111111111101, 27'b111111111111111111111111111, 27'b111111111111111110001011101, 27'b111111111111111111111111111, 27'b000000000000000000000000010, 27'b000000000000000000000000000, 27'b111111111111111111111010110, 27'b000000000000000000000010001, 27'b000000000000000001010110111, 27'b000000000000000000010011101, 27'b111111111111111111111111111, 27'b000000000000000000000000001, 27'b000000000000000000000111010, 27'b000000000000000000100111010, 27'b111111111111111101111000110, 27'b000000000000000001000101100, 27'b000000000000000011111110100, 27'b111111111111111111111111111, 27'b000000000000000000000110010, 27'b000000000000000000110010110, 27'b000000000000000001000111000}, 
{27'b000000000000000001100010100, 27'b000000000000000000000000000, 27'b111111111111111110010110011, 27'b111111111111111011111111001, 27'b111111111111110011010010111, 27'b000000000000000010001000010, 27'b000000000000000000000000011, 27'b111111111111110010110000110, 27'b000000000000000000100101001, 27'b111111111111111111111111101, 27'b000000000000000000000011110, 27'b111111111111111111111110010, 27'b000000000000000000001010110, 27'b000000000000000000000000001, 27'b111111111111111111101100101, 27'b111111111111111001111001001, 27'b111111111111111111111111111, 27'b000000000000000011100001001, 27'b000000000000000010000001011, 27'b000000000000000011000011110, 27'b111111111111111000111101110, 27'b111111111111111010010011100, 27'b000000000000000001111010111, 27'b111111111111111111011100010, 27'b111111111111111111010000110, 27'b000000000000000101101111001, 27'b111111111111111110011101000, 27'b111111111111111111111111101, 27'b111111111111111111111111110, 27'b000000000000000011011000001, 27'b111111111111111111111111110, 27'b000000000000000000000110011}, 
{27'b111111111111111100110101111, 27'b111111111111111000000111001, 27'b000000000000000000000000000, 27'b111111111111111111111101110, 27'b000000000000000101010100000, 27'b111111111111111011101100010, 27'b111111111111111100011101010, 27'b000000000000000001110110101, 27'b111111111111111111111111011, 27'b000000000000000010011000010, 27'b000000000000000001001011110, 27'b111111111111111110110010100, 27'b000000000000000000000000010, 27'b000000000000000000001110011, 27'b111111111111111111101010010, 27'b111111111111111011111100111, 27'b000000000000000010110011101, 27'b000000000000000000011101001, 27'b000000000000000100110000011, 27'b000000000000000001011000100, 27'b000000000000000000000000000, 27'b111111111111111111011001010, 27'b000000000000000010000001000, 27'b111111111111111110100111100, 27'b111111111111111011000100100, 27'b111111111111111111111001001, 27'b000000000000000010111101011, 27'b111111111111111111111111110, 27'b000000000000000000001000101, 27'b111111111111111110011111000, 27'b000000000000000010001100110, 27'b000000000000000100011010111}, 
{27'b000000000000000000001111100, 27'b000000000000000000000000001, 27'b000000000000000011100000100, 27'b000000000000000000001000100, 27'b111111111111111111010110010, 27'b000000000000000010111000110, 27'b000000000000000001011110011, 27'b111111111111111111111111101, 27'b000000000000000000000000110, 27'b111111111111111101110000011, 27'b111111111111111111001000000, 27'b111111111111111101010100101, 27'b111111111111111111111111110, 27'b000000000000000000110011101, 27'b111111111111111110111001011, 27'b000000000000001101011111011, 27'b000000000000000000000000010, 27'b111111111111111110011111101, 27'b111111111111111100111110110, 27'b111111111111111111110010011, 27'b000000000000000011001011011, 27'b000000000000000010000011000, 27'b000000000000000000000000001, 27'b111111111111111111111101011, 27'b000000000000000011100000110, 27'b000000000000000100010010100, 27'b000000000000000111111011001, 27'b000000000000000000001010100, 27'b000000000000000000000000001, 27'b000000000000000000000000011, 27'b111111111111111111110011110, 27'b111111111111111110110110110}, 
{27'b111111111111111101100000000, 27'b000000000000000000110001100, 27'b000000000000000000101000010, 27'b111111111111111100000010110, 27'b111111111111111011101100000, 27'b000000000000000111100000001, 27'b000000000000000000110010010, 27'b000000000000000000000000000, 27'b111111111111111101011011011, 27'b111111111111111110100101100, 27'b000000000000000010000100101, 27'b000000000000000001001000100, 27'b000000000000000000000000100, 27'b111111111111111110101111101, 27'b000000000000000100100100111, 27'b111111111111111111111111110, 27'b111111111111111111110010000, 27'b000000000000000000000000001, 27'b000000000000000000001101011, 27'b111111111111111111010000011, 27'b000000000000000001010000001, 27'b000000000000000000010000001, 27'b000000000000000001110100110, 27'b111111111111111111111111101, 27'b000000000000000000000011011, 27'b000000000000001010100001111, 27'b111111111111111111000110010, 27'b111111111111111111101000011, 27'b111111111111111111111111110, 27'b111111111111111110010000001, 27'b111111111111111111010110111, 27'b000000000000000010110100001}, 
{27'b000000000000000000111100010, 27'b000000000000000001001011111, 27'b000000000000000101001110010, 27'b111111111111111111010111010, 27'b000000000000000001100111011, 27'b000000000000000101100111010, 27'b000000000000000000000000101, 27'b111111111111111111100001111, 27'b000000000000000001111000110, 27'b111111111111111110001011011, 27'b111111111111111111111111111, 27'b111111111111111110000101111, 27'b000000000000000000000000010, 27'b000000000000000110010010101, 27'b111111111111111111101101111, 27'b000000000000000000000001101, 27'b000000000000000011110001110, 27'b000000000000000000000000101, 27'b000000000000000000000011000, 27'b111111111111111010111111101, 27'b111111111111111100000100100, 27'b111111111111111111011011000, 27'b111111111111111111111111111, 27'b111111111111111101101010100, 27'b111111111111111111011011000, 27'b111111111111111110101011100, 27'b111111111111111100110110111, 27'b111111111111111100100110011, 27'b000000000000000000011110110, 27'b000000000000000001110010010, 27'b111111111111111001101001001, 27'b000000000000000000000011010}, 
{27'b111111111111111011001110010, 27'b000000000000000000000000000, 27'b111111111111111111110000110, 27'b111111111111111111001101001, 27'b111111111111111111111111110, 27'b000000000000000010001000100, 27'b111111111111111110110000110, 27'b000000000000000100010101100, 27'b111111111111111010001100001, 27'b111111111111111111111111011, 27'b000000000000000000000000000, 27'b111111111111111111111111111, 27'b000000000000000000000000010, 27'b000000000000000000000000001, 27'b111111111111111111111100001, 27'b111111111111111110100011001, 27'b000000000000000001010001001, 27'b000000000000000010111011101, 27'b111111111111111111110110011, 27'b111111111111111011111110101, 27'b111111111111111111000011110, 27'b000000000000000001110010100, 27'b000000000000000001000000100, 27'b000000000000000000000000011, 27'b000000000000000000000011000, 27'b000000000000000001010011101, 27'b111111111111111100001010110, 27'b000000000000000000000000000, 27'b111111111111111111111111111, 27'b000000000000000000000011011, 27'b000000000000000000000000100, 27'b111111111111111101111111001}, 
{27'b111111111111111010100111110, 27'b111111111111111111111010000, 27'b111111111111111111111100111, 27'b111111111111111111101110001, 27'b111111111111111111111011000, 27'b000000000000000001101100000, 27'b000000000000000000000110110, 27'b000000000000000000100011011, 27'b000000000000000000100111000, 27'b000000000000000001000000011, 27'b000000000000000001010000110, 27'b000000000000000010100101000, 27'b000000000000000000011011011, 27'b111111111111111110011100111, 27'b000000000000000000000000100, 27'b000000000000000110000110100, 27'b000000000000000000000000010, 27'b000000000000000000000001001, 27'b111111111111111111111101011, 27'b000000000000000001110000101, 27'b000000000000000010010001110, 27'b000000000000000000011111100, 27'b000000000000000000101010001, 27'b111111111111111111100001100, 27'b111111111111111111011111000, 27'b000000000000000000011011001, 27'b111111111111111110111011010, 27'b111111111111111101111110010, 27'b000000000000000011010110100, 27'b111111111111111111100000100, 27'b000000000000000000100000011, 27'b111111111111111100111111101}, 
{27'b000000000000000000000000001, 27'b111111111111111111111111111, 27'b000000000000000000100110100, 27'b000000000000000000000000001, 27'b000000000000001110100000011, 27'b111111111111111111111111001, 27'b000000000000000000000000000, 27'b111111111111111111111111111, 27'b000000000000000001110000010, 27'b111111111111111110110011000, 27'b000000000000000000000000000, 27'b000000000000000000000000000, 27'b000000000000000000000001001, 27'b000000000000000010000100001, 27'b000000000000000000000000000, 27'b111111111111111101101011001, 27'b111111111111111111111111111, 27'b111111111111111110111011011, 27'b000000000000000101001111010, 27'b000000000000000000000000001, 27'b111111111111111111111111111, 27'b111111111111111111111111101, 27'b000000000000000000000000000, 27'b111111111111111111111111111, 27'b000000000000000000000000000, 27'b000000000000000001000101111, 27'b000000000000000000000000000, 27'b000000000000000000000000000, 27'b111111111111111111111111111, 27'b111111111111111111111111110, 27'b000000000000000000000000001, 27'b000000000000000000101010011}, 
{27'b111111111111111111111100100, 27'b000000000000000000011101101, 27'b111111111111111111111111001, 27'b000000000000000000110001000, 27'b111111111111111111010010100, 27'b111111111111111110000101110, 27'b111111111111111111000000000, 27'b000000000000000100011100011, 27'b000000000000000000000000010, 27'b000000000000000001100011001, 27'b111111111111111111110100101, 27'b000000000000000001000010011, 27'b111111111111111111011110000, 27'b111111111111111101011110101, 27'b111111111111111100111100111, 27'b000000000000000000001101011, 27'b111111111111111111111111111, 27'b111111111111111111011100010, 27'b000000000000000000000000000, 27'b000000000000000000000000011, 27'b111111111111111111111111011, 27'b000000000000000001001101100, 27'b000000000000000000100100100, 27'b111111111111111101111111001, 27'b000000000000000001110010011, 27'b111111111111111101010111100, 27'b000000000000000000000010001, 27'b000000000000000000000000000, 27'b111111111111111101010100010, 27'b000000000000000000000000000, 27'b000000000000000000101110101, 27'b111111111111111111100000001}, 
{27'b111111111111111111110100001, 27'b111111111111111110011010101, 27'b000000000000000000000000001, 27'b111111111111111111000010110, 27'b000000000000000011011101001, 27'b111111111111111111111111101, 27'b111111111111111111101010101, 27'b000000000000000001101101010, 27'b111111111111111001101111110, 27'b000000000000000000000000001, 27'b111111111111111111011000100, 27'b111111111111111111111101110, 27'b000000000000000101100111111, 27'b000000000000000011101010111, 27'b111111111111111110011010010, 27'b111111111111111111101010101, 27'b111111111111111111111111101, 27'b000000000000000000000000101, 27'b111111111111111111111111110, 27'b000000000000000000000000010, 27'b000000000000000000000000001, 27'b111111111111111101110100111, 27'b111111111111111110000110001, 27'b000000000000000010000110000, 27'b000000000000000000000000000, 27'b111111111111111101110011101, 27'b000000000000000000011001000, 27'b111111111111111110101101101, 27'b111111111111111111011101111, 27'b000000000000000010001011001, 27'b000000000000000000000000100, 27'b111111111111111100000010111}, 
{27'b000000000000001010001001111, 27'b000000000000000101011110001, 27'b111111111111111100000000101, 27'b000000000000000000000011010, 27'b111111111111111010011101101, 27'b000000000000000000000000000, 27'b000000000000000011100100001, 27'b000000000000000000011111110, 27'b000000000000000011100101001, 27'b111111111111111111111111101, 27'b111111111111111101100001011, 27'b111111111111111110101111100, 27'b000000000000000010010001001, 27'b000000000000000000011100010, 27'b111111111111111110011011011, 27'b000000000000000010000110111, 27'b000000000000001000100100000, 27'b111111111111111101111010110, 27'b111111111111111011010000110, 27'b000000000000000000000000000, 27'b111111111111111111100010101, 27'b111111111111111101001011001, 27'b111111111111111111110011100, 27'b111111111111111111111110011, 27'b000000000000000001011000000, 27'b111111111111111010001110111, 27'b000000000000000001011011000, 27'b111111111111111111111110111, 27'b000000000000000000000000010, 27'b000000000000000001101111101, 27'b111111111111111111100010011, 27'b000000000000000000111101000}, 
{27'b111111111111111110100001001, 27'b111111111111111100111011011, 27'b111111111111111111011010110, 27'b111111111111111101010100101, 27'b111111111111111111101110011, 27'b000000000000000000110010011, 27'b000000000000000000000000001, 27'b111111111111111111110100011, 27'b000000000000000000100110100, 27'b111111111111111111111100011, 27'b000000000000000000000000001, 27'b111111111111111100100001110, 27'b000000000000000001101000011, 27'b000000000000000001010010010, 27'b111111111111111110010111001, 27'b000000000000000111000110001, 27'b111111111111111111111111110, 27'b000000000000000000000000001, 27'b111111111111111111111011111, 27'b000000000000000000000000000, 27'b000000000000000101000011101, 27'b111111111111111000011110000, 27'b111111111111111110010001000, 27'b111111111111111111000110101, 27'b111111111111111111101100111, 27'b000000000000000011001001110, 27'b111111111111111111001010010, 27'b000000000000000000010010000, 27'b000000000000000111101111111, 27'b111111111111110111110011001, 27'b111111111111111010001000000, 27'b000000000000000000010110111}, 
{27'b000000000000000000010001001, 27'b111111111111111111000011110, 27'b111111111111111111111111111, 27'b000000000000000000000000001, 27'b111111111111110100011111110, 27'b111111111111110110010011000, 27'b000000000000000000000001100, 27'b111111111111111111111111110, 27'b111111111111111011110000100, 27'b000000000000000000011001010, 27'b000000000000000000000000000, 27'b111111111111111111100011110, 27'b000000000000000000000000000, 27'b111111111111111111000100001, 27'b111111111111111111001010001, 27'b111111111111111110111001011, 27'b111111111111111101101001011, 27'b000000000000000100100001000, 27'b000000000000000000000000000, 27'b000000000000000000101111010, 27'b111111111111111111111111100, 27'b111111111111111110110111110, 27'b000000000000000000000000000, 27'b111111111111111110100111001, 27'b000000000000000011100000110, 27'b111111111111110110000010101, 27'b000000000000000011100001011, 27'b111111111111111111111111111, 27'b111111111111111111111011000, 27'b000000000000000011001100110, 27'b111111111111111111111111111, 27'b000000000000000011110001111}, 
{27'b111111111111111111111111110, 27'b000000000000000000000101010, 27'b111111111111111111010011110, 27'b000000000000000001001100111, 27'b000000000000000000111000101, 27'b111111111111111010100001110, 27'b000000000000000000000000001, 27'b000000000000000001000001111, 27'b000000000000001001010001100, 27'b111111111111111111110110110, 27'b000000000000000000000000000, 27'b000000000000000000111001101, 27'b000000000000000101101111100, 27'b111111111111111111011111011, 27'b000000000000000000001110010, 27'b000000000000000001100111011, 27'b111111111111111111111111111, 27'b000000000000000000011100011, 27'b111111111111111111111111101, 27'b000000000000000000000000111, 27'b111111111111111011100111101, 27'b000000000000000000100111010, 27'b000000000000000001000111111, 27'b000000000000000000010111010, 27'b111111111111111111111111110, 27'b000000000000000011011111100, 27'b000000000000000000000100100, 27'b000000000000000010000001000, 27'b111111111111111001010100011, 27'b000000000000000001101001010, 27'b000000000000000110010101001, 27'b000000000000000000000101110}, 
{27'b111111111111111010011000101, 27'b000000000000000011011000001, 27'b111111111111111011110101010, 27'b000000000000000001111101111, 27'b111111111111111110010100000, 27'b000000000000000000000000010, 27'b000000000000000111111101100, 27'b111111111111111100010001101, 27'b111111111111111011010101110, 27'b000000000000000010101111011, 27'b111111111111111100011011111, 27'b111111111111111111100111111, 27'b111111111111111111111111000, 27'b000000000000000101100000010, 27'b111111111111111111111110011, 27'b111111111111111011001011000, 27'b111111111111111111111111111, 27'b000000000000000111000011011, 27'b111111111111111000011101101, 27'b111111111111111111100111001, 27'b000000000000000101000100001, 27'b111111111111111010001100101, 27'b000000000000000000110110010, 27'b111111111111111111110000100, 27'b000000000000000100010101111, 27'b111111111111110111110111001, 27'b111111111111111010001100100, 27'b111111111111111100110111001, 27'b111111111111111111111111111, 27'b000000000000000001101010000, 27'b000000000000000000011001101, 27'b000000000000000010110110101}, 
{27'b111111111111111110100011000, 27'b000000000000000000110101001, 27'b111111111111111111111111110, 27'b000000000000000010011001011, 27'b111111111111111111011001001, 27'b000000000000000011101000011, 27'b000000000000000000000010000, 27'b111111111111111111110100100, 27'b111111111111111111111101111, 27'b000000000000000000000001001, 27'b000000000000000000000000000, 27'b111111111111111111111111111, 27'b111111111111111111111110000, 27'b000000000000001000010100101, 27'b000000000000000000001100111, 27'b000000000000000011000001011, 27'b000000000000000000000000010, 27'b111111111111111100100111010, 27'b111111111111111110110001110, 27'b111111111111111111111111111, 27'b111111111111111111101111000, 27'b000000000000000000101011001, 27'b111111111111111111111111111, 27'b111111111111111101000010010, 27'b111111111111111111111111111, 27'b000000000000000100101110101, 27'b000000000000000100111101101, 27'b111111111111111111111111111, 27'b111111111111111111101111010, 27'b000000000000000000000000000, 27'b111111111111111111111111011, 27'b111111111111111110011101010}, 
{27'b111111111111111110101101010, 27'b000000000000000000000000000, 27'b000000000000000100010111100, 27'b000000000000000000000000000, 27'b000000000000000000000000000, 27'b111111111111111110001011101, 27'b000000000000000000000000010, 27'b111111111111110010001011100, 27'b000000000000000011011100101, 27'b000000000000000000001110000, 27'b000000000000000000011011010, 27'b111111111111111010001111100, 27'b000000000000000000000011011, 27'b111111111111111101110011010, 27'b111111111111111111011110000, 27'b000000000000000000000000001, 27'b000000000000000000010100000, 27'b000000000000000000000000001, 27'b000000000000000001110011000, 27'b000000000000000000000000010, 27'b111111111111111111110110111, 27'b000000000000000101010001001, 27'b000000000000000110000001100, 27'b111111111111111100011101110, 27'b111111111111111101101110100, 27'b000000000000000011111111100, 27'b111111111111111011000111000, 27'b000000000000000000011110000, 27'b111111111111111111111111011, 27'b111111111111111111111111111, 27'b111111111111111111111111110, 27'b000000000000000010111100100}, 
{27'b111111111111111110001011110, 27'b111111111111111111111111011, 27'b111111111111111100001011000, 27'b111111111111111100110001001, 27'b111111111111111111110001111, 27'b111111111111111101110101111, 27'b000000000000000000000000000, 27'b000000000000000001011101010, 27'b111111111111111100001010100, 27'b111111111111111110101010101, 27'b111111111111111111001101001, 27'b000000000000000000000000010, 27'b000000000000000000011100100, 27'b111111111111111111110101111, 27'b111111111111111111000001100, 27'b000000000000000001100001111, 27'b000000000000000011100100001, 27'b000000000000000010000110010, 27'b111111111111111101111010000, 27'b000000000000000000110001111, 27'b111111111111111111110011111, 27'b111111111111111111100010110, 27'b000000000000000000010111000, 27'b000000000000000000010000010, 27'b111111111111111110111000111, 27'b000000000000000001011011001, 27'b111111111111111110100011001, 27'b000000000000000000111101010, 27'b111111111111111111111111110, 27'b111111111111111011010001101, 27'b111111111111111111100101000, 27'b000000000000000011100110010}, 
{27'b111111111111111111100100011, 27'b111111111111111110101011010, 27'b000000000000000001001110110, 27'b000000000000000100000011001, 27'b000000000000000001010110110, 27'b000000000000000001010100010, 27'b000000000000000000101111110, 27'b111111111111111100110001101, 27'b111111111111111100101101111, 27'b000000000000000001000110000, 27'b000000000000000000001100011, 27'b000000000000000000101100001, 27'b000000000000000000010110110, 27'b000000000000000000000101100, 27'b000000000000000011010010000, 27'b000000000000000000000111100, 27'b111111111111111111001000110, 27'b000000000000000001101001110, 27'b111111111111111111100001101, 27'b111111111111111111011011011, 27'b000000000000000001110000101, 27'b111111111111111110000001000, 27'b111111111111111111100100101, 27'b000000000000000010000010000, 27'b000000000000000000010110101, 27'b111111111111111110010010110, 27'b111111111111111100110101011, 27'b111111111111111111110011111, 27'b111111111111111011100010001, 27'b000000000000000000111101100, 27'b000000000000000001101000001, 27'b000000000000000000000001001}, 
{27'b111111111111111111110010000, 27'b111111111111111111101011110, 27'b111111111111111111110011110, 27'b111111111111111111011100100, 27'b111111111111111101111001010, 27'b111111111111111101110000010, 27'b000000000000000001000000101, 27'b000000000000000000001000011, 27'b111111111111111101000101001, 27'b000000000000000010101011011, 27'b111111111111111111101010101, 27'b111111111111111111111111011, 27'b111111111111111110001111001, 27'b000000000000000000000101010, 27'b000000000000000000011110001, 27'b111111111111111111001010001, 27'b111111111111111111101111101, 27'b111111111111111111010101010, 27'b111111111111111110101101101, 27'b000000000000000000000000010, 27'b111111111111111101110000001, 27'b000000000000000001101000010, 27'b111111111111111100100111011, 27'b000000000000000000000101000, 27'b000000000000000000101010111, 27'b000000000000000001111110111, 27'b000000000000000000011011001, 27'b000000000000000000000110001, 27'b000000000000000100101011000, 27'b000000000000000000110100110, 27'b000000000000000000000000010, 27'b000000000000000001010101110}, 
{27'b111111111111111111101100001, 27'b000000000000000100000010110, 27'b111111111111111111111111111, 27'b111111111111111111011110010, 27'b111111111111111100100101001, 27'b111111111111111110110011000, 27'b000000000000000110100101010, 27'b111111111111110100111110010, 27'b111111111111111010011010000, 27'b111111111111111100110011101, 27'b111111111111111100011111010, 27'b111111111111111011111100011, 27'b111111111111111111111111011, 27'b000000000000000111101111111, 27'b111111111111111111100101001, 27'b000000000000000000000000000, 27'b111111111111111100100111110, 27'b000000000000000111001000011, 27'b111111111111111001011001010, 27'b000000000000000000000000001, 27'b111111111111111111111111101, 27'b111111111111111010100111101, 27'b000000000000000000000000001, 27'b111111111111111111111111111, 27'b000000000000000000111001100, 27'b111111111111111111000101001, 27'b111111111111111101101000101, 27'b111111111111111111111111111, 27'b000000000000000010110010110, 27'b000000000000000000000011011, 27'b111111111111111110101101110, 27'b000000000000000000000000110}, 
{27'b000000000000000101111000110, 27'b111111111111111110001101011, 27'b000000000000000010000111000, 27'b111111111111111111011110111, 27'b000000000000000001001110000, 27'b111111111111111111111100001, 27'b111111111111111111111101000, 27'b111111111111111110100000110, 27'b000000000000000000000000010, 27'b000000000000000001011110011, 27'b111111111111111111111111111, 27'b111111111111111111000011111, 27'b111111111111111111111111100, 27'b000000000000000011101010001, 27'b000000000000000000010011101, 27'b000000000000000000101001011, 27'b000000000000000000011000100, 27'b111111111111111111100111011, 27'b000000000000000000010100110, 27'b000000000000000000000000001, 27'b111111111111111111110110110, 27'b111111111111111111111111111, 27'b111111111111111011000111000, 27'b111111111111111111111111111, 27'b000000000000000000111011001, 27'b111111111111111110001000111, 27'b111111111111111101110101100, 27'b111111111111111111111111111, 27'b111111111111111111111111001, 27'b000000000000001000111011001, 27'b111111111111111011011011011, 27'b111111111111111110001001000}, 
{27'b111111111111111111010010111, 27'b111111111111111110010110010, 27'b111111111111111110111101111, 27'b000000000000000000100101001, 27'b000000000000000010001110110, 27'b111111111111111101111011000, 27'b111111111111111111111110101, 27'b111111111111111100011110111, 27'b000000000000000000111110001, 27'b000000000000000010001011010, 27'b111111111111111100100101011, 27'b111111111111111011111101001, 27'b000000000000000000011000011, 27'b111111111111110101000100001, 27'b111111111111111110110010110, 27'b111111111111111110000001100, 27'b111111111111111100110101011, 27'b111111111111111111111111101, 27'b000000000000000010001001011, 27'b000000000000000000000000000, 27'b111111111111111111010001010, 27'b111111111111111111010010010, 27'b000000000000000000000000000, 27'b000000000000000000000000000, 27'b111111111111111111000011100, 27'b111111111111110011111011100, 27'b111111111111110111000111010, 27'b111111111111111011101000111, 27'b000000000000000000111001010, 27'b000000000000000011010011001, 27'b111111111111111111111111101, 27'b000000000000000011110110000}, 
{27'b111111111111111110100001101, 27'b111111111111111100100100000, 27'b000000000000000010100111101, 27'b000000000000000001001100011, 27'b000000000000000000101100011, 27'b111111111111111110100001110, 27'b111111111111111111011110100, 27'b000000000000000001100100111, 27'b000000000000001000100111111, 27'b111111111111111101010000101, 27'b111111111111111111111111111, 27'b111111111111111111111111111, 27'b000000000000000001111000011, 27'b111111111111111111000111110, 27'b111111111111111111101101101, 27'b111111111111111111101110111, 27'b111111111111111110011001101, 27'b111111111111111111111111000, 27'b000000000000000000000000000, 27'b000000000000000011101000000, 27'b111111111111111101110111110, 27'b111111111111111111111100111, 27'b000000000000000010000011101, 27'b111111111111111111110101100, 27'b000000000000000000000000000, 27'b000000000000001000011010111, 27'b000000000000000101001100000, 27'b000000000000000000000011010, 27'b000000000000000000000000010, 27'b111111111111111001010001000, 27'b111111111111111110111010000, 27'b111111111111111111111111111}, 
{27'b000000000000000000001111011, 27'b000000000000000000110001011, 27'b111111111111111111110001111, 27'b000000000000000000000000000, 27'b000000000000000011101100111, 27'b111111111111111000010001001, 27'b000000000000000000000000001, 27'b111111111111111110011110101, 27'b000000000000000010111110111, 27'b000000000000000000000000000, 27'b111111111111111111101101000, 27'b000000000000000000000000000, 27'b000000000000000000000000010, 27'b111111111111111111111111110, 27'b000000000000000000000101111, 27'b111111111111111110010001111, 27'b000000000000000100001001101, 27'b111111111111111111111010011, 27'b111111111111111111110000001, 27'b111111111111111111111111111, 27'b000000000000000000000000010, 27'b111111111111111111111000001, 27'b000000000000000000000000010, 27'b111111111111111111111111111, 27'b000000000000000000001101001, 27'b111111111111111010111011011, 27'b000000000000000000110100111, 27'b000000000000000010111011101, 27'b111111111111111111111100101, 27'b000000000000000001100000100, 27'b111111111111111111111111101, 27'b000000000000000001001100100}, 
{27'b111111111111111100110001111, 27'b000000000000000000001001010, 27'b111111111111111000010010000, 27'b000000000000000000000111000, 27'b111111111111111111001100110, 27'b111111111111111111010111010, 27'b111111111111111111111110101, 27'b111111111111111110100010101, 27'b111111111111111111011011001, 27'b111111111111111110111101000, 27'b000000000000000000110000001, 27'b000000000000000000011011100, 27'b111111111111111101001010011, 27'b000000000000000000000000100, 27'b111111111111111111111110000, 27'b111111111111111111110111101, 27'b000000000000000001001000001, 27'b111111111111111111101011010, 27'b111111111111111111100011110, 27'b111111111111111111100010010, 27'b111111111111111111111111001, 27'b000000000000000100010101100, 27'b111111111111111111111111111, 27'b000000000000000000000000000, 27'b111111111111111111110110011, 27'b000000000000000101000100111, 27'b000000000000000011000001001, 27'b000000000000000000100010110, 27'b111111111111111110011101010, 27'b111111111111111111110101110, 27'b000000000000000001000010110, 27'b000000000000000000111010111}, 
{27'b000000000000000000100010111, 27'b000000000000000000101000000, 27'b111111111111111111111111110, 27'b000000000000000000000000011, 27'b111111111111111000100000000, 27'b000000000000000000101100101, 27'b000000000000000000011001011, 27'b111111111111111111111111101, 27'b000000000000000000000000101, 27'b111111111111111101010010011, 27'b111111111111111111111111111, 27'b000000000000000000000000000, 27'b111111111111111101011011010, 27'b000000000000000000000000001, 27'b000000000000000000000000010, 27'b000000000000000000000000010, 27'b000000000000000000000000000, 27'b111111111111111010010011101, 27'b000000000000000000001001110, 27'b111111111111111111111111011, 27'b111111111111111111111111100, 27'b000000000000000000000000001, 27'b000000000000000010000100000, 27'b111111111111111111111111111, 27'b000000000000000000000000001, 27'b000000000000000111010010110, 27'b000000000000000101011100010, 27'b000000000000000000000000001, 27'b000000000000000000000000001, 27'b111111111111111100010000110, 27'b000000000000000000000000011, 27'b111111111111111111111111111}, 
{27'b000000000000000001001101100, 27'b000000000000000000110110000, 27'b000000000000000100000011001, 27'b111111111111111100000001110, 27'b000000000000000010000111100, 27'b000000000000000001111001100, 27'b000000000000000000000110011, 27'b000000000000000011000100011, 27'b000000000000000000001100001, 27'b111111111111111111110011101, 27'b000000000000000000100110001, 27'b000000000000000000000101111, 27'b111111111111111111111111011, 27'b000000000000000001111011100, 27'b111111111111111111111010010, 27'b111111111111111111010111011, 27'b000000000000000000000000101, 27'b000000000000000000100000100, 27'b111111111111111111001110101, 27'b000000000000000001100101000, 27'b000000000000000000100001010, 27'b111111111111110110101101101, 27'b111111111111111110001010110, 27'b000000000000000001011101100, 27'b111111111111111111111111111, 27'b111111111111110111111010111, 27'b111111111111111101111110110, 27'b111111111111111111101000011, 27'b111111111111111111111111010, 27'b111111111111111111000101100, 27'b000000000000000000000000000, 27'b111111111111111111010111011}, 
{27'b000000000000000000000001111, 27'b111111111111111111111111111, 27'b111111111111111110100010010, 27'b111111111111111101010011101, 27'b000000000000000000101010111, 27'b000000000000000000000000001, 27'b000000000000000001100001100, 27'b111111111111111111111010001, 27'b000000000000000011111111100, 27'b111111111111111111111011111, 27'b000000000000000000000000000, 27'b111111111111111010100000010, 27'b111111111111111111111111100, 27'b000000000000000010000000111, 27'b111111111111111111111111110, 27'b111111111111111011110101000, 27'b000000000000000000000000000, 27'b111111111111111111110100011, 27'b000000000000000100001101001, 27'b111111111111111111111111111, 27'b111111111111111001000000111, 27'b111111111111111111111111111, 27'b000000000000000100001000001, 27'b111111111111111111111111111, 27'b111111111111111111111111111, 27'b000000000000000010001110001, 27'b111111111111111110011111111, 27'b000000000000000001000110110, 27'b000000000000000000000000001, 27'b111111111111111100110001101, 27'b000000000000000000000000000, 27'b000000000000000000000010100}, 
{27'b111111111111111100100010100, 27'b000000000000000000000001001, 27'b000000000000000000000000100, 27'b111111111111111111111001110, 27'b000000000000000111111011101, 27'b111111111111111110000000110, 27'b111111111111111111111010010, 27'b111111111111111111111000100, 27'b111111111111111111010010001, 27'b111111111111111111001100011, 27'b000000000000000001000010110, 27'b000000000000000010001000000, 27'b111111111111111111011010010, 27'b000000000000000011111111100, 27'b000000000000000000000000001, 27'b111111111111111111111111100, 27'b111111111111111011011101000, 27'b111111111111111111111111011, 27'b000000000000000000000000011, 27'b111111111111111110101110011, 27'b000000000000000000000010001, 27'b000000000000000000100110001, 27'b000000000000000000001101101, 27'b111111111111111111110110101, 27'b111111111111111111001011111, 27'b111111111111111100110000010, 27'b111111111111111011010001000, 27'b000000000000000000000000010, 27'b111111111111111110001100000, 27'b000000000000000000101000110, 27'b111111111111111111111111101, 27'b000000000000000001001101011}, 
{27'b111111111111111001011000111, 27'b111111111111111101011111110, 27'b111111111111111101100000000, 27'b000000000000000000000000000, 27'b000000000000001001001000111, 27'b111111111111111100011100000, 27'b000000000000000000000000000, 27'b111111111111111111001000100, 27'b111111111111111001011100010, 27'b000000000000000010001101110, 27'b111111111111111111111111111, 27'b000000000000001001000100110, 27'b000000000000000000000000011, 27'b111111111111111111001111011, 27'b111111111111111111111111101, 27'b000000000000000000100000011, 27'b111111111111111111101100111, 27'b000000000000000000000000011, 27'b111111111111111111010000010, 27'b000000000000000111111011010, 27'b000000000000000000100111101, 27'b111111111111111111010101010, 27'b000000000000000001110000001, 27'b111111111111111111111111101, 27'b111111111111111111111111111, 27'b111111111111111110011100011, 27'b111111111111111111010000000, 27'b111111111111111000100000111, 27'b111111111111111101101100001, 27'b111111111111111111111111111, 27'b111111111111111111111110111, 27'b111111111111111111000011111}, 
{27'b000000000000000011100111010, 27'b111111111111110011001101010, 27'b111111111111110100011010001, 27'b111111111111111101010001110, 27'b000000000000001010101101011, 27'b111111111111111111111111111, 27'b111111111111111010011101000, 27'b000000000000000100001111001, 27'b000000000000000000111100110, 27'b000000000000000000000000111, 27'b000000000000000011010101011, 27'b111111111111111011101010000, 27'b000000000000000000000000111, 27'b000000000000000000000100011, 27'b111111111111111111011111111, 27'b000000000000000000010010011, 27'b111111111111111110010101101, 27'b111111111111110001010000011, 27'b000000000000000010101011110, 27'b000000000000000101100001001, 27'b000000000000000100001111011, 27'b000000000000000000000010101, 27'b000000000000000000011101110, 27'b111111111111111001100011011, 27'b111111111111110101111000000, 27'b111111111111111111111010111, 27'b111111111111111011001101000, 27'b111111111111111000101011001, 27'b111111111111111100111000011, 27'b111111111111110001111101111, 27'b000000000000000110101101010, 27'b000000000000000110110111100}, 
{27'b000000000000000000000000010, 27'b000000000000000000000000101, 27'b000000000000000000000010010, 27'b000000000000000000000000001, 27'b000000000000000100001001001, 27'b111111111111111101000000100, 27'b000000000000000000010010001, 27'b000000000000000001001010101, 27'b111111111111111010011010101, 27'b000000000000000000100101100, 27'b111111111111111111111011011, 27'b111111111111111111111111000, 27'b111111111111111111111111110, 27'b000000000000000011110101010, 27'b000000000000000000110101001, 27'b000000000000000000010110010, 27'b000000000000000000111111010, 27'b000000000000000101010101010, 27'b111111111111111100100000010, 27'b000000000000000000000000000, 27'b111111111111111101010111110, 27'b111111111111111111111111101, 27'b000000000000000101000010001, 27'b000000000000000000001000010, 27'b111111111111111111111101000, 27'b111111111111110111000001011, 27'b111111111111111111110110100, 27'b111111111111111101100001111, 27'b111111111111111111000001100, 27'b000000000000000000000011101, 27'b000000000000000010001010010, 27'b000000000000000001101010001}, 
{27'b111111111111111111010011101, 27'b000000000000000010001001001, 27'b111111111111111011001000111, 27'b000000000000000000010101001, 27'b000000000000000011000110010, 27'b111111111111111111010111100, 27'b111111111111111111111011010, 27'b000000000000000010100111001, 27'b000000000000000000000000010, 27'b111111111111111111111111110, 27'b111111111111111110111101000, 27'b000000000000000000000000000, 27'b000000000000000000000000011, 27'b111111111111111111011100111, 27'b111111111111111110000011011, 27'b111111111111111110111100000, 27'b111111111111111111000110010, 27'b111111111111111110111111101, 27'b111111111111111110001111100, 27'b000000000000000000000000000, 27'b111111111111111111111111101, 27'b111111111111111111010010001, 27'b111111111111111110111011110, 27'b000000000000000110010111010, 27'b000000000000000000000000000, 27'b111111111111111010001111011, 27'b111111111111111111110111010, 27'b000000000000000001111110001, 27'b000000000000000000000000011, 27'b000000000000000000000000000, 27'b000000000000000100000000111, 27'b111111111111111111111111100}, 
{27'b111111111111111111111111111, 27'b000000000000000000000100001, 27'b111111111111111111111111101, 27'b111111111111111101100000000, 27'b111111111111110010001111000, 27'b000000000000000000000000111, 27'b000000000000000000000000010, 27'b111111111111111111111001010, 27'b111111111111110110011010000, 27'b000000000000000001010011100, 27'b111111111111111110011011100, 27'b111111111111111111111111111, 27'b000000000000000000000000011, 27'b111111111111111010000101001, 27'b111111111111111111010001000, 27'b111111111111111111111111101, 27'b000000000000000000000001011, 27'b000000000000000000001000011, 27'b000000000000000000100101001, 27'b000000000000000101100001100, 27'b111111111111111110000101100, 27'b111111111111111011001101110, 27'b000000000000000000000000000, 27'b111111111111111011110111111, 27'b111111111111111110011010111, 27'b111111111111111100010011000, 27'b111111111111111111111000011, 27'b111111111111111111110011001, 27'b111111111111111111101101011, 27'b111111111111111000011101100, 27'b111111111111111111011101000, 27'b000000000000000011111000000}, 
{27'b000000000000000001110011111, 27'b000000000000000011100000011, 27'b111111111111111111111101111, 27'b000000000000000010100011001, 27'b111111111111111100101000000, 27'b111111111111111110000000100, 27'b000000000000000001100001111, 27'b000000000000000001000110010, 27'b111111111111111111001111110, 27'b111111111111111111111111111, 27'b111111111111111111111111111, 27'b111111111111111111111111110, 27'b111111111111111111111111101, 27'b111111111111111010110111111, 27'b111111111111111111111111111, 27'b000000000000000010010011101, 27'b111111111111111110001010111, 27'b000000000000000000100011101, 27'b111111111111111111111110101, 27'b111111111111111111111110111, 27'b000000000000000011010100011, 27'b111111111111111010110001000, 27'b000000000000000100011111100, 27'b000000000000000000110000101, 27'b000000000000000000000000010, 27'b000000000000000011011000111, 27'b000000000000000000000011001, 27'b111111111111111111011011000, 27'b111111111111111001111010010, 27'b111111111111111110001111111, 27'b111111111111111101010001101, 27'b000000000000000010110101110}, 
{27'b000000000000000000000000000, 27'b000000000000000000000111011, 27'b111111111111111010001001010, 27'b111111111111111111111101100, 27'b000000000000000011010011101, 27'b111111111111111101101111000, 27'b111111111111111111110011101, 27'b111111111111111111111111111, 27'b000000000000000000010100110, 27'b000000000000000000000000000, 27'b000000000000000000000000000, 27'b111111111111111100101111010, 27'b000000000000000001100010010, 27'b000000000000000000000110001, 27'b000000000000000000000000001, 27'b000000000000000000100110010, 27'b111111111111111111111111101, 27'b111111111111111101100111101, 27'b000000000000000000010010010, 27'b000000000000000000000000001, 27'b111111111111111111011100110, 27'b111111111111111111101001100, 27'b000000000000000100101111011, 27'b111111111111111111111111111, 27'b000000000000000000000000000, 27'b111111111111111011010100010, 27'b111111111111111010110001010, 27'b000000000000000011110111001, 27'b111111111111111111111110101, 27'b111111111111111111111111101, 27'b000000000000000000011100010, 27'b000000000000000100100001011}, 
{27'b111111111111111010100011000, 27'b111111111111111111111111111, 27'b111111111111111100100110001, 27'b000000000000000000000100011, 27'b111111111111111010010110001, 27'b000000000000000000000000000, 27'b111111111111111111111111101, 27'b111111111111111110111101000, 27'b111111111111110111011110111, 27'b111111111111111111100101101, 27'b000000000000000000000000000, 27'b111111111111111111110111100, 27'b111111111111111111111111101, 27'b000000000000000000000000000, 27'b111111111111111111110111001, 27'b111111111111111111001101000, 27'b111111111111111101101000111, 27'b111111111111111110011110010, 27'b000000000000000001000011110, 27'b111111111111111111111101100, 27'b111111111111111111100110000, 27'b000000000000000000000000000, 27'b000000000000000101011000110, 27'b111111111111111111111111110, 27'b000000000000000010011001000, 27'b000000000000000001011101111, 27'b111111111111111101110011000, 27'b000000000000000011011010011, 27'b111111111111111111010001001, 27'b000000000000000000000000000, 27'b111111111111111111111110110, 27'b000000000000001001010100000}, 
{27'b111111111111111010111110011, 27'b000000000000000000011110011, 27'b000000000000000000110011111, 27'b111111111111111111100011010, 27'b000000000000000011111010000, 27'b111111111111111011001010100, 27'b111111111111111111111000110, 27'b000000000000000100001111111, 27'b000000000000000010100011001, 27'b000000000000000000001001011, 27'b111111111111111111111111111, 27'b111111111111111110111001111, 27'b111111111111111110100100011, 27'b111111111111111110111101110, 27'b111111111111111111001101001, 27'b000000000000000001011100011, 27'b111111111111111111111111111, 27'b000000000000000000001000010, 27'b000000000000000010010000101, 27'b000000000000000000000000000, 27'b000000000000000000000000000, 27'b000000000000000000001111010, 27'b000000000000000100000010000, 27'b000000000000000000101110110, 27'b000000000000000000000110110, 27'b111111111111111110010001110, 27'b111111111111111111111111111, 27'b000000000000000000000000000, 27'b111111111111111111110001100, 27'b111111111111111111110011101, 27'b111111111111111111111111101, 27'b000000000000000001000101001}, 
{27'b111111111111111111111111110, 27'b000000000000000000000011111, 27'b111111111111111100100110111, 27'b111111111111111110110011101, 27'b000000000000000100100000111, 27'b111111111111111111111111101, 27'b111111111111111110110000101, 27'b000000000000000011111010010, 27'b111111111111111111001001110, 27'b000000000000000100101010101, 27'b000000000000000001010111100, 27'b111111111111111110000100111, 27'b000000000000000000000000100, 27'b000000000000000000000011100, 27'b111111111111111111110000111, 27'b000000000000000000010101110, 27'b111111111111111110110001000, 27'b111111111111111011110010011, 27'b000000000000000100011100100, 27'b000000000000000010011111000, 27'b000000000000001010001001111, 27'b000000000000000011001101100, 27'b000000000000000011111110000, 27'b111111111111111111111111110, 27'b000000000000000000000000000, 27'b000000000000000000000000000, 27'b000000000000000000111010101, 27'b000000000000000001010001001, 27'b111111111111111001010001111, 27'b111111111111111111111111110, 27'b111111111111111111111010110, 27'b111111111111111111111001010}, 
{27'b000000000000000000000000100, 27'b111111111111111110100110010, 27'b111111111111111110010101111, 27'b000000000000000000000000000, 27'b111111111111111100000110100, 27'b000000000000000000000000000, 27'b000000000000000011000100000, 27'b000000000000000001101111110, 27'b000000000000000000110110011, 27'b111111111111111110011010111, 27'b000000000000000000000000000, 27'b111111111111111111111111111, 27'b111111111111111111111111110, 27'b111111111111111111111111110, 27'b111111111111111111010100010, 27'b000000000000000011001110111, 27'b111111111111111111111111111, 27'b111111111111111111111111011, 27'b111111111111111011001010011, 27'b000000000000000000000000001, 27'b111111111111111100111010111, 27'b111111111111111111111110111, 27'b000000000000000000000000001, 27'b111111111111111111111011110, 27'b000000000000000000001111011, 27'b000000000000000000010001110, 27'b000000000000000000011100100, 27'b000000000000000010001101101, 27'b111111111111111110111101011, 27'b111111111111111111111000001, 27'b111111111111111000110100100, 27'b000000000000000001010000101}, 
{27'b000000000000000111000100011, 27'b111111111111111111110111000, 27'b000000000000000001000011110, 27'b111111111111111110010100110, 27'b111111111111111110101000100, 27'b000000000000000000100010001, 27'b000000000000000010100100000, 27'b000000000000000000000000000, 27'b000000000000001000011011101, 27'b000000000000000000000000010, 27'b111111111111111111101010000, 27'b000000000000000000010011010, 27'b000000000000000001100000010, 27'b111111111111111111111101010, 27'b000000000000000000110110100, 27'b000000000000000001101001110, 27'b111111111111111111111011100, 27'b111111111111111000111000001, 27'b111111111111111111000110010, 27'b111111111111111111111110010, 27'b000000000000000001110111000, 27'b000000000000000000000001101, 27'b111111111111111111111111100, 27'b000000000000000001110011001, 27'b000000000000000000010010011, 27'b111111111111111011110010000, 27'b111111111111111110010110110, 27'b000000000000000010000111011, 27'b111111111111111111100011000, 27'b000000000000000100001000010, 27'b111111111111111111111110111, 27'b111111111111111101001000111}, 
{27'b000000000000000000001101010, 27'b000000000000000001101000010, 27'b111111111111111111111111111, 27'b111111111111111111011000010, 27'b111111111111111010010110100, 27'b111111111111111111111111100, 27'b000000000000000000101111001, 27'b111111111111111111010000110, 27'b000000000000000010101000110, 27'b111111111111111111011101000, 27'b111111111111111111111111001, 27'b111111111111111111011101110, 27'b111111111111111111111111110, 27'b111111111111111111011010000, 27'b000000000000000000000000000, 27'b000000000000000101000000100, 27'b000000000000000000000000000, 27'b111111111111111111111110001, 27'b111111111111111111111111110, 27'b111111111111111111111111110, 27'b111111111111111111111111110, 27'b111111111111111111111111100, 27'b000000000000000000100010111, 27'b000000000000000010000000111, 27'b000000000000000000000000000, 27'b000000000000000000000100010, 27'b000000000000000000100001001, 27'b111111111111111111111111011, 27'b000000000000000000000000000, 27'b000000000000000000010100111, 27'b000000000000000000000001100, 27'b000000000000000001100011001}, 
{27'b111111111111111011000011110, 27'b000000000000000010000101011, 27'b000000000000000000010010011, 27'b111111111111111110010100011, 27'b111111111111111001100111001, 27'b111111111111111111101101010, 27'b000000000000000001000100100, 27'b111111111111111001101001000, 27'b000000000000001000001011110, 27'b000000000000000001001001011, 27'b000000000000000000010000000, 27'b000000000000000001100000100, 27'b000000000000000000101101011, 27'b000000000000000000000000101, 27'b000000000000000110100001100, 27'b111111111111111110101001110, 27'b000000000000000000000101010, 27'b000000000000000000000000000, 27'b111111111111111111111001001, 27'b000000000000000000000011110, 27'b111111111111111001000101111, 27'b000000000000000000010001010, 27'b000000000000000010011100100, 27'b000000000000000000100110011, 27'b000000000000000000100100111, 27'b111111111111110101011111111, 27'b111111111111111010100010111, 27'b111111111111111100001001100, 27'b000000000000000000000010101, 27'b111111111111111111111110001, 27'b000000000000000101001101101, 27'b111111111111111100101110010}, 
{27'b111111111111111111110010110, 27'b111111111111111100111000111, 27'b111111111111111110010110001, 27'b111111111111111001011101100, 27'b111111111111111011110101100, 27'b000000000000000101011000010, 27'b000000000000000100111101010, 27'b111111111111111101010001110, 27'b000000000000000000101010100, 27'b111111111111111111011000010, 27'b111111111111111110011111110, 27'b111111111111111011111110100, 27'b000000000000000001101001100, 27'b111111111111111011011101000, 27'b000000000000000011000001010, 27'b111111111111111111111111101, 27'b000000000000000101010111111, 27'b111111111111111111111111111, 27'b111111111111111111111000000, 27'b111111111111111101110101011, 27'b111111111111111111010101011, 27'b111111111111111110111101111, 27'b111111111111111011101111111, 27'b000000000000000001010100010, 27'b111111111111111111111111111, 27'b111111111111111111111001100, 27'b111111111111111100010110010, 27'b000000000000000101000010011, 27'b000000000000000100011101110, 27'b111111111111111110100011011, 27'b111111111111110101111010010, 27'b000000000000000010010010010}, 
{27'b000000000000000000000000011, 27'b111111111111111111100101110, 27'b111111111111111111111111110, 27'b111111111111111110011100011, 27'b000000000000000000011101001, 27'b000000000000000000001001010, 27'b000000000000000001000111010, 27'b000000000000000000000101111, 27'b000000000000000001111000101, 27'b111111111111111111111111000, 27'b000000000000000000000000000, 27'b000000000000000001100001101, 27'b000000000000000000000001111, 27'b000000000000000000001100100, 27'b111111111111111101111000011, 27'b111111111111111110010001101, 27'b000000000000000000000000000, 27'b000000000000000010111010000, 27'b000000000000000000111010001, 27'b000000000000000010000000110, 27'b111111111111111111101111000, 27'b111111111111111101011100010, 27'b111111111111111111111111110, 27'b000000000000000001001100000, 27'b111111111111111111111111110, 27'b000000000000000000100001001, 27'b111111111111111111111011000, 27'b000000000000000001000101001, 27'b000000000000000000000000001, 27'b000000000000000001010101001, 27'b111111111111111001111011011, 27'b111111111111111111111111111}, 
{27'b000000000000000100111101110, 27'b111111111111111111110110110, 27'b000000000000000010011001100, 27'b111111111111111011000111011, 27'b111111111111111100111010010, 27'b111111111111111111111111111, 27'b111111111111111111111111110, 27'b000000000000000000011100000, 27'b000000000000000000000010011, 27'b111111111111111101111111000, 27'b000000000000000000000000000, 27'b000000000000000000000010000, 27'b000000000000000000000000000, 27'b000000000000000000000000010, 27'b111111111111111101111011110, 27'b000000000000000010010010000, 27'b111111111111111111111110010, 27'b111111111111111111100000010, 27'b000000000000000000000000001, 27'b000000000000000001111010111, 27'b111111111111111100110010011, 27'b000000000000000001110110111, 27'b000000000000000010001111011, 27'b000000000000000010000100000, 27'b111111111111111111111111111, 27'b000000000000001000110100101, 27'b111111111111111101100011001, 27'b000000000000000101110100001, 27'b111111111111111111001011001, 27'b111111111111111010001110101, 27'b111111111111111101001110011, 27'b000000000000000010001110110}, 
{27'b111111111111110111010011110, 27'b111111111111111111100100101, 27'b111111111111111101100010010, 27'b111111111111111111111111111, 27'b000000000000000100001011000, 27'b111111111111111101001001001, 27'b111111111111111111000010101, 27'b000000000000000011110011111, 27'b000000000000000001100000110, 27'b111111111111111100001100010, 27'b000000000000000000000000001, 27'b111111111111111111100011001, 27'b111111111111111111110101111, 27'b000000000000000010001100110, 27'b111111111111111100000100011, 27'b111111111111111111110100100, 27'b000000000000000000000000000, 27'b111111111111111111111111010, 27'b111111111111111111101111100, 27'b000000000000000000000000000, 27'b111111111111111100111101010, 27'b111111111111111111111111110, 27'b000000000000000000000000000, 27'b111111111111111010101111110, 27'b000000000000000001000111111, 27'b000000000000001001111010101, 27'b000000000000000101100010001, 27'b111111111111111111011011010, 27'b111111111111111101011011100, 27'b111111111111111000110100100, 27'b000000000000000000000000010, 27'b111111111111111111001110000}, 
{27'b000000000000000000010101111, 27'b000000000000000011011010110, 27'b000000000000000000010101110, 27'b111111111111111101100101010, 27'b000000000000000000000100101, 27'b111111111111111111100101111, 27'b000000000000000000000000001, 27'b000000000000000011010101011, 27'b000000000000000011011100000, 27'b111111111111111101110111001, 27'b000000000000000010001111110, 27'b000000000000000000011000100, 27'b111111111111111111111111111, 27'b111111111111111111110001011, 27'b111111111111111101011101011, 27'b000000000000000100000011000, 27'b111111111111111111010100100, 27'b111111111111111010110101001, 27'b000000000000000001110101000, 27'b111111111111111111111111110, 27'b111111111111111111111111110, 27'b000000000000000001110111101, 27'b111111111111111110110011111, 27'b111111111111111111111011000, 27'b111111111111111111001011001, 27'b000000000000000001011010010, 27'b111111111111111101110000010, 27'b000000000000000010001001010, 27'b111111111111111010001011100, 27'b000000000000000001010010011, 27'b111111111111111111111111100, 27'b000000000000000010100000011}, 
{27'b111111111111111111010100000, 27'b000000000000000000000000100, 27'b000000000000000001011011001, 27'b000000000000000000000000000, 27'b111111111111111111000001100, 27'b111111111111111111111101000, 27'b000000000000000001101001000, 27'b111111111111111111111111111, 27'b000000000000000000000000001, 27'b000000000000000000000101001, 27'b000000000000000000000000001, 27'b000000000000000000010100011, 27'b111111111111111110010011001, 27'b000000000000000000001010101, 27'b000000000000000001110001011, 27'b000000000000000000101111110, 27'b000000000000000001101100000, 27'b111111111111111111111111011, 27'b111111111111111111111110101, 27'b000000000000000010000011000, 27'b000000000000000011111101010, 27'b111111111111111110011011110, 27'b000000000000000000000000000, 27'b111111111111111111111101111, 27'b000000000000000000001011101, 27'b111111111111111000100111111, 27'b111111111111111111111111001, 27'b111111111111111110110111100, 27'b111111111111111111111111110, 27'b000000000000001001000010001, 27'b000000000000000000000000010, 27'b111111111111111100101101001}, 
{27'b111111111111111111100100100, 27'b111111111111111110000101110, 27'b111111111111111111110110111, 27'b000000000000000000000111001, 27'b000000000000000001011100111, 27'b111111111111111111111111111, 27'b000000000000000000000000001, 27'b111111111111111111101000010, 27'b000000000000000001001000010, 27'b111111111111111111110111100, 27'b000000000000000000000000001, 27'b000000000000000000100000011, 27'b000000000000000100101110000, 27'b111111111111111110010111100, 27'b000000000000000000001100111, 27'b111111111111110010011011011, 27'b111111111111111111110100100, 27'b111111111111111111000010000, 27'b000000000000000000001000001, 27'b111111111111111111001100111, 27'b000000000000000001011110001, 27'b111111111111111100011010100, 27'b000000000000000001110100111, 27'b000000000000000001101011111, 27'b111111111111111111110010100, 27'b111111111111110100100111111, 27'b111111111111111100010101111, 27'b111111111111111111101001101, 27'b111111111111111111101101001, 27'b000000000000000110001111111, 27'b111111111111111111111010000, 27'b000000000000000010011101110}, 
{27'b000000000000000000110000000, 27'b000000000000000000000000001, 27'b000000000000000010110010010, 27'b111111111111111110001011110, 27'b111111111111111110111001100, 27'b000000000000000011110011100, 27'b111111111111111101011100010, 27'b000000000000000000111010111, 27'b111111111111111011000011001, 27'b000000000000000000001000111, 27'b000000000000000000010001001, 27'b111111111111111110101010000, 27'b000000000000000000000000100, 27'b000000000000000000000000000, 27'b111111111111111100111111101, 27'b000000000000000110111010110, 27'b111111111111111100000011010, 27'b111111111111111111110011110, 27'b000000000000000001111001101, 27'b111111111111111111111111110, 27'b000000000000000001000110111, 27'b111111111111111000010101011, 27'b000000000000000101000000101, 27'b111111111111111111111111111, 27'b111111111111111110000001001, 27'b000000000000000111110000010, 27'b000000000000000010010101100, 27'b111111111111111101011110011, 27'b111111111111111101110110010, 27'b111111111111110111011001111, 27'b111111111111111111110101100, 27'b000000000000000000010000010}, 
{27'b111111111111111111111111111, 27'b000000000000000000000110101, 27'b111111111111111111011100011, 27'b111111111111111011101101100, 27'b111111111111111111111111101, 27'b111111111111111001101110001, 27'b000000000000000000000000010, 27'b000000000000000100110110111, 27'b000000000000000011111010001, 27'b000000000000000000010011010, 27'b000000000000000000000000000, 27'b111111111111111110001111001, 27'b000000000000000101010100000, 27'b111111111111111111111111111, 27'b111111111111111111111111101, 27'b111111111111111111111111100, 27'b000000000000000110111100010, 27'b000000000000000000000001101, 27'b111111111111111111010111010, 27'b111111111111111111001011101, 27'b111111111111111010110110011, 27'b000000000000000010000110110, 27'b000000000000000000000000000, 27'b000000000000000000000000000, 27'b000000000000000000100000011, 27'b111111111111111110110111001, 27'b111111111111111000101000010, 27'b000000000000000100011010100, 27'b111111111111111000111001111, 27'b000000000000000000110100010, 27'b111111111111111110101111001, 27'b000000000000000000000000000}, 
{27'b000000000000000000111110110, 27'b000000000000000010111110111, 27'b000000000000000000001001111, 27'b111111111111111111111100111, 27'b111111111111111000101001101, 27'b000000000000000000000000111, 27'b111111111111111111111111111, 27'b000000000000000011111000000, 27'b000000000000000100011011101, 27'b111111111111111111111111110, 27'b111111111111111111111111110, 27'b111111111111111111111110101, 27'b000000000000000000000000001, 27'b000000000000000000000010000, 27'b000000000000000000000000000, 27'b000000000000000000000000001, 27'b000000000000000000000000011, 27'b111111111111111111111111010, 27'b000000000000000010101110000, 27'b111111111111111110010110100, 27'b111111111111111001000101101, 27'b111111111111111111011110000, 27'b111111111111111110011010110, 27'b111111111111111110011111111, 27'b111111111111111110111001000, 27'b111111111111111111111111000, 27'b111111111111111110111111100, 27'b111111111111111111101001100, 27'b111111111111111111110101010, 27'b000000000000000010010000110, 27'b111111111111111111111111101, 27'b000000000000000111011010100}
};

localparam logic signed [26:0] bias [32] = '{
27'b000000000000010111100101101,  // 1.474280834197998
27'b000000000000001011000100000,  // 0.6914801001548767
27'b000000000000010111000011001,  // 1.4406442642211914
27'b000000000000010110100001110,  // 1.408045768737793
27'b000000000000001111110010001,  // 0.9864811301231384
27'b000000000000001101110100010,  // 0.8636202812194824
27'b111111111111110110001001110,  // -0.6153604388237
27'b000000000000000111101111100,  // 0.4839226007461548
27'b000000000000000111110001111,  // 0.4862793982028961
27'b000000000000000101111100100,  // 0.37162142992019653
27'b000000000000000111010110111,  // 0.45989668369293213
27'b000000000000010100110011000,  // 1.2998151779174805
27'b111111111111101111101111000,  // -1.016528844833374
27'b111111111111111010010111000,  // -0.35249894857406616
27'b000000000000000111001000100,  // 0.44582197070121765
27'b111111111111111110001101010,  // -0.1119980737566948
27'b111111111111111110111011001,  // -0.06717441976070404
27'b000000000000000000000100111,  // 0.00487547367811203
27'b000000000000000011000111010,  // 0.1946917623281479
27'b111111111111110011100001100,  // -0.7796769738197327
27'b000000000000001011101010001,  // 0.7287401556968689
27'b000000000000011011011100000,  // 1.714877724647522
27'b111111111111100110011100100,  // -1.5971007347106934
27'b000000000000000001001011101,  // 0.07393483817577362
27'b000000000000000101001010010,  // 0.3225609362125397
27'b000000000000001101100001100,  // 0.8453295230865479
27'b000000000000001110011000001,  // 0.898597240447998
27'b000000000000000100000100111,  // 0.2548799514770508
27'b000000000000001111100100111,  // 0.9735668301582336
27'b000000000000010010000001001,  // 1.1261906623840332
27'b000000000000000111001010011,  // 0.44768181443214417
27'b111111111111011010000111100   // -2.3676068782806396
};
endpackage