// Width: 8
// NFRAC: 4
package dense_1_8_4;

localparam logic signed [7:0] weights [16][64] = '{ 
{8'b00000100, 8'b11110101, 8'b11111101, 8'b11111100, 8'b11111001, 8'b00000001, 8'b11101111, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000000, 8'b11111001, 8'b11111111, 8'b00000011, 8'b00000000, 8'b11111011, 8'b00000011, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000110, 8'b11111010, 8'b11111111, 8'b00000111, 8'b11111010, 8'b11110101, 8'b11111011, 8'b11111100, 8'b11111110, 8'b11111111, 8'b00000000, 8'b00000011, 8'b00000011, 8'b11111111, 8'b00000000, 8'b00000100, 8'b11111111, 8'b11111011, 8'b00000000, 8'b00000011, 8'b11111111, 8'b00000100, 8'b11111011, 8'b00001110, 8'b11111111, 8'b00000111, 8'b00000000, 8'b00000010, 8'b00000011, 8'b11111111, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000001, 8'b11111110, 8'b11111011, 8'b00001000, 8'b11111000, 8'b00000111, 8'b11111010, 8'b00001100, 8'b11111111, 8'b00000000, 8'b00000001}, 
{8'b00000000, 8'b11111010, 8'b11111101, 8'b11111011, 8'b11111010, 8'b00000001, 8'b11110011, 8'b11111111, 8'b11111100, 8'b00000010, 8'b00000000, 8'b11111110, 8'b00000011, 8'b00000000, 8'b11111111, 8'b00000011, 8'b11111111, 8'b00000000, 8'b11111101, 8'b11111011, 8'b00000111, 8'b11111110, 8'b00000000, 8'b00001011, 8'b00000100, 8'b11111100, 8'b11111100, 8'b11111111, 8'b11111110, 8'b11111001, 8'b11111111, 8'b00000111, 8'b00000100, 8'b00001000, 8'b00001010, 8'b00000000, 8'b11111110, 8'b11111001, 8'b00000000, 8'b00000011, 8'b00000000, 8'b00000011, 8'b11111100, 8'b00000100, 8'b00000010, 8'b00000000, 8'b11111010, 8'b00000001, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00010010, 8'b11111110, 8'b11111110, 8'b11111111, 8'b11111111, 8'b00000100, 8'b11111010, 8'b00001111, 8'b00000000, 8'b00001000, 8'b00000011, 8'b00001101, 8'b00000010}, 
{8'b11111111, 8'b00000000, 8'b11111110, 8'b11111101, 8'b11111101, 8'b00000000, 8'b00010111, 8'b11111111, 8'b11101011, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111100, 8'b00000000, 8'b11111111, 8'b00000010, 8'b00001110, 8'b11111111, 8'b00000001, 8'b00000000, 8'b00000110, 8'b11110100, 8'b00001001, 8'b11110100, 8'b00001111, 8'b11111010, 8'b11111100, 8'b11110100, 8'b00010100, 8'b00000100, 8'b00000000, 8'b00001000, 8'b00010000, 8'b11101100, 8'b11111110, 8'b00000000, 8'b11111100, 8'b00001110, 8'b11111111, 8'b00000101, 8'b00000101, 8'b00000101, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000010, 8'b11111011, 8'b11111101, 8'b11111111, 8'b00000110, 8'b11111101, 8'b00000010, 8'b11111111, 8'b00000010, 8'b11111101, 8'b11111111, 8'b11111011, 8'b11110101, 8'b11111111, 8'b00000000, 8'b00011000, 8'b00000000, 8'b11111111, 8'b11111011}, 
{8'b11111000, 8'b11111010, 8'b11110100, 8'b00000100, 8'b11111010, 8'b11101010, 8'b11111110, 8'b11111011, 8'b00000011, 8'b11111111, 8'b00010100, 8'b11111110, 8'b11110011, 8'b00001001, 8'b00000000, 8'b11111111, 8'b11111000, 8'b11111111, 8'b00000000, 8'b11111100, 8'b11101101, 8'b11111110, 8'b11110100, 8'b00000011, 8'b11111001, 8'b11110001, 8'b00000101, 8'b00001011, 8'b00010100, 8'b11111000, 8'b11110110, 8'b00000001, 8'b00001000, 8'b11110010, 8'b11111010, 8'b00000000, 8'b11110100, 8'b00000011, 8'b11111000, 8'b00000001, 8'b00000111, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00001000, 8'b11111100, 8'b11111111, 8'b11111010, 8'b11111111, 8'b11111110, 8'b11110110, 8'b00000001, 8'b11111111, 8'b00000011, 8'b00000101, 8'b00001010, 8'b11110000, 8'b11110001, 8'b11110100, 8'b00001101, 8'b00011011, 8'b11110001, 8'b11111111, 8'b00000110}, 
{8'b00000101, 8'b11110110, 8'b11111011, 8'b11111111, 8'b11111101, 8'b00000101, 8'b00000011, 8'b11111111, 8'b11110110, 8'b11111100, 8'b11111010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000101, 8'b00000010, 8'b11111001, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11111110, 8'b00000001, 8'b11111111, 8'b00010001, 8'b11111101, 8'b11111011, 8'b11111001, 8'b00000000, 8'b00000010, 8'b00000001, 8'b00000100, 8'b11111111, 8'b00000001, 8'b00000010, 8'b11111111, 8'b00000000, 8'b00001110, 8'b11111011, 8'b11111110, 8'b00000110, 8'b00000011, 8'b11111000, 8'b00000000, 8'b11101110, 8'b11111111, 8'b11111110, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000011, 8'b11111111, 8'b00000101, 8'b11111100, 8'b11110100, 8'b11111000, 8'b11110111, 8'b11110110, 8'b00001011, 8'b00010101, 8'b00001100, 8'b00000001, 8'b11111111}, 
{8'b11111000, 8'b11110101, 8'b00000000, 8'b00000100, 8'b00000100, 8'b11111100, 8'b00001001, 8'b11111111, 8'b00000011, 8'b11111111, 8'b11111111, 8'b11111110, 8'b11111101, 8'b00001001, 8'b11111110, 8'b00000000, 8'b11110110, 8'b11111010, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111010, 8'b11111010, 8'b00000111, 8'b11111010, 8'b11111111, 8'b00000100, 8'b11111110, 8'b11110001, 8'b11111111, 8'b11111110, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000000, 8'b11111110, 8'b11111011, 8'b11111111, 8'b11111101, 8'b11110111, 8'b00000110, 8'b00000000, 8'b00001001, 8'b00000000, 8'b11111111, 8'b00000001, 8'b11111001, 8'b00000011, 8'b00000000, 8'b11111110, 8'b11111010, 8'b00000110, 8'b11111111, 8'b00000101, 8'b00000011, 8'b00000011, 8'b11111111, 8'b11111111, 8'b11110011, 8'b11111101, 8'b11111111, 8'b11111111}, 
{8'b11111011, 8'b11111010, 8'b11111001, 8'b11111110, 8'b11111101, 8'b00000001, 8'b11110100, 8'b11111101, 8'b11111100, 8'b11111111, 8'b11111011, 8'b00000101, 8'b00000000, 8'b00000010, 8'b00000100, 8'b00000000, 8'b00001100, 8'b00000001, 8'b00000011, 8'b00000100, 8'b11111101, 8'b00000101, 8'b11111100, 8'b11110111, 8'b00000010, 8'b00001000, 8'b11111111, 8'b00000000, 8'b11110000, 8'b00000100, 8'b00000100, 8'b11111010, 8'b00000111, 8'b00001010, 8'b00000000, 8'b00000101, 8'b11111111, 8'b00000100, 8'b00000011, 8'b00000000, 8'b11111110, 8'b11111010, 8'b00000010, 8'b00000111, 8'b00001000, 8'b11111101, 8'b11111110, 8'b11111100, 8'b11111101, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b11111101, 8'b00001100, 8'b00000101, 8'b11111111, 8'b00000110, 8'b00000011, 8'b11100101, 8'b11110110, 8'b11111101, 8'b11111111}, 
{8'b00000000, 8'b00000011, 8'b11111111, 8'b11111111, 8'b11111010, 8'b11111111, 8'b11111011, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b11111001, 8'b11111110, 8'b00000000, 8'b11111111, 8'b11111000, 8'b11110010, 8'b11111111, 8'b11110110, 8'b11111000, 8'b11111001, 8'b00000101, 8'b00000000, 8'b11111101, 8'b11111001, 8'b00000010, 8'b00000000, 8'b00000111, 8'b00001100, 8'b11111111, 8'b00000000, 8'b00000011, 8'b11110101, 8'b11111010, 8'b00000000, 8'b00000001, 8'b11111011, 8'b00000011, 8'b00000010, 8'b11111101, 8'b11111001, 8'b11111111, 8'b00000000, 8'b11111101, 8'b00000000, 8'b00000011, 8'b11111110, 8'b00000000, 8'b00000000, 8'b11111100, 8'b11111001, 8'b00000110, 8'b00000010, 8'b11111101, 8'b00000010, 8'b11111111, 8'b11111000, 8'b11111101, 8'b11111111, 8'b11111110, 8'b00001101, 8'b00000011, 8'b11111111, 8'b11111111}, 
{8'b00000000, 8'b00001001, 8'b11110110, 8'b11111100, 8'b00000101, 8'b11111100, 8'b00010011, 8'b11111011, 8'b11111111, 8'b00000100, 8'b00000100, 8'b11111111, 8'b11111111, 8'b11111000, 8'b00000100, 8'b00000010, 8'b11111100, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000100, 8'b11111000, 8'b00000110, 8'b00001001, 8'b11111110, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00001011, 8'b00000000, 8'b11111011, 8'b00000000, 8'b00000110, 8'b11110011, 8'b11110111, 8'b00000011, 8'b00000010, 8'b11110110, 8'b11111100, 8'b11111100, 8'b00000110, 8'b00000110, 8'b00000000, 8'b11111011, 8'b00000000, 8'b00000110, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000011, 8'b11111111, 8'b11111100, 8'b00000101, 8'b11111100, 8'b00000100, 8'b00001001, 8'b00000000, 8'b00000100, 8'b11111001, 8'b11111010, 8'b00001101, 8'b11111101, 8'b00000000, 8'b11111110}, 
{8'b00000000, 8'b11111000, 8'b00000101, 8'b11111011, 8'b11111111, 8'b00000011, 8'b11110110, 8'b00000011, 8'b00000111, 8'b00000010, 8'b00000101, 8'b00000101, 8'b11111011, 8'b11111110, 8'b11111111, 8'b00000000, 8'b11110000, 8'b00000101, 8'b11111111, 8'b00000000, 8'b11111010, 8'b00000001, 8'b00000010, 8'b11111111, 8'b11111000, 8'b11111111, 8'b11111110, 8'b00010011, 8'b11110101, 8'b00000001, 8'b00000001, 8'b11111111, 8'b11111100, 8'b00000001, 8'b11111110, 8'b11111101, 8'b11111101, 8'b11111100, 8'b11111111, 8'b11111011, 8'b00000101, 8'b00000001, 8'b00000111, 8'b00000001, 8'b00000000, 8'b11111011, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000011, 8'b00000010, 8'b00000100, 8'b11111111, 8'b11111011, 8'b00000000, 8'b00000000, 8'b00000101, 8'b11111100, 8'b11110111, 8'b00001000, 8'b11111011, 8'b00010010, 8'b11111111, 8'b11111010}, 
{8'b11110110, 8'b11111111, 8'b11111001, 8'b00000011, 8'b00000100, 8'b11111110, 8'b00001000, 8'b11111101, 8'b11111000, 8'b11111010, 8'b11111011, 8'b11111000, 8'b11111100, 8'b00000011, 8'b00000000, 8'b00000000, 8'b00001101, 8'b11111111, 8'b11111111, 8'b00000110, 8'b00000100, 8'b11110110, 8'b11111001, 8'b00000011, 8'b11111001, 8'b11111111, 8'b11111011, 8'b11111010, 8'b11111001, 8'b00000100, 8'b00000011, 8'b11111101, 8'b11111110, 8'b11110000, 8'b11111101, 8'b00000000, 8'b11111101, 8'b11111011, 8'b11111111, 8'b00000001, 8'b11111110, 8'b11111111, 8'b11111111, 8'b11110101, 8'b00000000, 8'b00000000, 8'b00000101, 8'b11111110, 8'b00000110, 8'b11111100, 8'b00000100, 8'b11111111, 8'b00000011, 8'b11111001, 8'b11111111, 8'b00001000, 8'b00000101, 8'b00000100, 8'b00000000, 8'b11111001, 8'b11111011, 8'b11110101, 8'b11111111, 8'b00000001}, 
{8'b00000100, 8'b00000000, 8'b00000010, 8'b11111111, 8'b00000010, 8'b11111101, 8'b00000011, 8'b00000000, 8'b00000010, 8'b00000101, 8'b11111011, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11110101, 8'b11111011, 8'b00001010, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111001, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000101, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111100, 8'b11110101, 8'b00000100, 8'b00000101, 8'b11111111, 8'b11111100, 8'b00000000, 8'b11110101, 8'b11111111, 8'b11111111, 8'b00000011, 8'b11111101, 8'b11111111, 8'b00001101, 8'b00000111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111100, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000110, 8'b00000101, 8'b00001010, 8'b11111101, 8'b00000110, 8'b00000010, 8'b11111010, 8'b00000001, 8'b11111001, 8'b11111000, 8'b11111000}, 
{8'b00000000, 8'b00000011, 8'b11111100, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11110101, 8'b11111111, 8'b00000100, 8'b00000011, 8'b00000011, 8'b11111001, 8'b11111110, 8'b00000100, 8'b11111111, 8'b00000000, 8'b11110010, 8'b11111111, 8'b00000101, 8'b00000001, 8'b00000011, 8'b11111110, 8'b00000011, 8'b00000110, 8'b11111010, 8'b11111011, 8'b11111111, 8'b11111110, 8'b00000001, 8'b00000000, 8'b11111111, 8'b00000101, 8'b11110100, 8'b00000101, 8'b00001000, 8'b00000001, 8'b00000001, 8'b11111110, 8'b00000001, 8'b11111110, 8'b11111011, 8'b11111111, 8'b00000010, 8'b00001011, 8'b11110010, 8'b11111000, 8'b00000011, 8'b11111110, 8'b00000111, 8'b11111100, 8'b11111010, 8'b11111011, 8'b11111111, 8'b00000001, 8'b11111101, 8'b11110010, 8'b11111101, 8'b11111111, 8'b00000000, 8'b11110110, 8'b00010001, 8'b11110111, 8'b00001000, 8'b00000010}, 
{8'b00000001, 8'b11111100, 8'b00001010, 8'b11111011, 8'b11111000, 8'b00000001, 8'b00000100, 8'b00000100, 8'b11111101, 8'b11111101, 8'b00000000, 8'b00000011, 8'b00000011, 8'b00000000, 8'b11111100, 8'b00000010, 8'b00000111, 8'b11111111, 8'b11111011, 8'b00000000, 8'b00000001, 8'b00000000, 8'b11111011, 8'b00000001, 8'b00001100, 8'b00000000, 8'b00000010, 8'b11110011, 8'b11111110, 8'b00000000, 8'b11111100, 8'b11111011, 8'b00000111, 8'b11111111, 8'b11111111, 8'b11111011, 8'b00000010, 8'b00000100, 8'b11111111, 8'b11111111, 8'b11111101, 8'b00000011, 8'b00000000, 8'b11110101, 8'b00000100, 8'b00000110, 8'b11111111, 8'b00000000, 8'b11111001, 8'b11111110, 8'b11111111, 8'b11111010, 8'b00000000, 8'b11111101, 8'b00000000, 8'b11110010, 8'b11111111, 8'b11111111, 8'b00000100, 8'b00001001, 8'b11110100, 8'b00001000, 8'b00000000, 8'b11111110}, 
{8'b00000100, 8'b00010011, 8'b00000111, 8'b00000100, 8'b11111000, 8'b11111010, 8'b11010110, 8'b11111000, 8'b00000110, 8'b11111111, 8'b00000100, 8'b00001101, 8'b00000001, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111100, 8'b11111100, 8'b00000011, 8'b11110111, 8'b11110101, 8'b11111110, 8'b11110110, 8'b00000000, 8'b11011011, 8'b00001101, 8'b00001111, 8'b00001001, 8'b11100100, 8'b11111010, 8'b11110100, 8'b11110010, 8'b11010111, 8'b00001010, 8'b11111111, 8'b00000101, 8'b00000000, 8'b11101001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00010000, 8'b11111100, 8'b11110101, 8'b00001110, 8'b11111000, 8'b11111010, 8'b11111001, 8'b00000111, 8'b00001000, 8'b11111110, 8'b11111010, 8'b11111111, 8'b11111110, 8'b00000000, 8'b11111001, 8'b00001001, 8'b00010001, 8'b00001011, 8'b11110001, 8'b11000100, 8'b00001110, 8'b00000001, 8'b00000101}, 
{8'b11111100, 8'b00000101, 8'b00000101, 8'b11111111, 8'b11111010, 8'b11111110, 8'b11111001, 8'b11111111, 8'b00000010, 8'b11111110, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111101, 8'b11111111, 8'b11111110, 8'b00000101, 8'b11111111, 8'b11110101, 8'b00000111, 8'b00001001, 8'b00000110, 8'b11111010, 8'b11111101, 8'b11111010, 8'b11111011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000101, 8'b00000000, 8'b00000110, 8'b11111111, 8'b00000000, 8'b00000100, 8'b00000010, 8'b11111110, 8'b11111111, 8'b00000000, 8'b11111011, 8'b11111100, 8'b11111110, 8'b11111010, 8'b00000111, 8'b00000000, 8'b11111111, 8'b11111110, 8'b11111101, 8'b11110011, 8'b11111111, 8'b11111100, 8'b11111101, 8'b11111110, 8'b00000100, 8'b00001010, 8'b00000010, 8'b11111111, 8'b11111010, 8'b11111111, 8'b00000000, 8'b00000101, 8'b11111111, 8'b00000000, 8'b00000000}
};

localparam logic signed [7:0] bias [64] = '{
8'b11111111,  // -0.037350185215473175
8'b00000100,  // 0.27355897426605225
8'b11111110,  // -0.12378914654254913
8'b11111110,  // -0.064457006752491
8'b00000000,  // 0.05452875792980194
8'b00000001,  // 0.11671770364046097
8'b00000010,  // 0.13640816509723663
8'b00000001,  // 0.07482525706291199
8'b00000000,  // 0.04674031585454941
8'b11111100,  // -0.20146161317825317
8'b11111110,  // -0.09910125285387039
8'b00000010,  // 0.15104414522647858
8'b11111110,  // -0.10221704095602036
8'b11111101,  // -0.1461549550294876
8'b11111110,  // -0.08641516417264938
8'b00000010,  // 0.16613510251045227
8'b11111110,  // -0.0836295336484909
8'b11111111,  // -0.05756539851427078
8'b11111111,  // -0.03229188174009323
8'b11111111,  // -0.028388574719429016
8'b00000010,  // 0.1260243058204651
8'b11111111,  // -0.037064336240291595
8'b00000011,  // 0.19336333870887756
8'b00000000,  // 0.02124214917421341
8'b00000111,  // 0.4985624849796295
8'b00000000,  // 0.0158411655575037
8'b11111110,  // -0.08296407759189606
8'b00000001,  // 0.11056788265705109
8'b00000000,  // 0.01173810102045536
8'b11111110,  // -0.10843746364116669
8'b00000100,  // 0.27439257502555847
8'b00000001,  // 0.09199801832437515
8'b00000100,  // 0.27419957518577576
8'b00000100,  // 0.27063727378845215
8'b11111100,  // -0.24828937649726868
8'b00000001,  // 0.07818280160427094
8'b11111111,  // -0.005749030504375696
8'b00000001,  // 0.10850494354963303
8'b00000010,  // 0.13591453433036804
8'b11111110,  // -0.12088628858327866
8'b11111111,  // -0.05666546896100044
8'b00000001,  // 0.09311636537313461
8'b00000000,  // 0.05477767437696457
8'b00000000,  // 0.029585206881165504
8'b11111011,  // -0.31209176778793335
8'b11111110,  // -0.08465463668107986
8'b11111101,  // -0.16775836050510406
8'b00000010,  // 0.14762157201766968
8'b11111100,  // -0.23618532717227936
8'b00000001,  // 0.06535740196704865
8'b11111101,  // -0.12853026390075684
8'b11111101,  // -0.13802281022071838
8'b11111101,  // -0.15156887471675873
8'b00000001,  // 0.07979883998632431
8'b00000010,  // 0.18141601979732513
8'b11111111,  // -0.054039113223552704
8'b11111111,  // -0.010052933357656002
8'b00000001,  // 0.06611225008964539
8'b00000000,  // 0.05053366720676422
8'b00000000,  // 0.026860840618610382
8'b00000000,  // 0.03283466026186943
8'b00000010,  // 0.15558314323425293
8'b11111011,  // -0.2863388657569885
8'b11111110   // -0.08769102394580841
};
endpackage