// Width: 19
// NFRAC: 9
package dense_2_19_9;

localparam logic signed [18:0] weights [64][32] = '{ 
{19'b0000000000010001001, 19'b0000000000000000100, 19'b1111111111110011110, 19'b1111111111111110101, 19'b0000000000010000101, 19'b0000000000000000000, 19'b1111111111110110110, 19'b1111111111111111111, 19'b1111111111101110011, 19'b0000000000000101000, 19'b0000000000000000000, 19'b1111111111111111101, 19'b1111111111111111111, 19'b1111111111110011001, 19'b1111111111111100110, 19'b1111111111101111001, 19'b0000000000000000000, 19'b1111111111111111001, 19'b1111111111110011110, 19'b1111111111110101110, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111111111011, 19'b1111111111111111110, 19'b0000000000000000000, 19'b0000000000000110011, 19'b0000000000011000101, 19'b0000000000001011001, 19'b1111111111111111111, 19'b0000000000000011001, 19'b1111111111100101110, 19'b0000000000000000000}, 
{19'b1111111111111001100, 19'b1111111111110110000, 19'b1111111111110111001, 19'b1111111111111100011, 19'b1111111111111111101, 19'b0000000000000010110, 19'b1111111111110001101, 19'b0000000000000000010, 19'b0000000000000000010, 19'b1111111111111011111, 19'b0000000000001001111, 19'b1111111111111101001, 19'b1111111111111100001, 19'b1111111111110010000, 19'b0000000000000000011, 19'b1111111111111100111, 19'b0000000000000000110, 19'b1111111111110011100, 19'b0000000000001010111, 19'b0000000000001110101, 19'b1111111111111101111, 19'b1111111111111111101, 19'b1111111111111111111, 19'b0000000000000001100, 19'b1111111111111011011, 19'b0000000000010001100, 19'b0000000000001111110, 19'b0000000000000000100, 19'b0000000000000001110, 19'b1111111111100000110, 19'b0000000000000000011, 19'b0000000000000000000}, 
{19'b0000000000000100101, 19'b1111111111111000101, 19'b1111111111110111101, 19'b1111111111111101010, 19'b1111111111111011000, 19'b1111111111111010100, 19'b1111111111110100001, 19'b0000000000000000010, 19'b1111111111110111010, 19'b0000000000000000100, 19'b0000000000000000001, 19'b1111111111111010110, 19'b0000000000000101110, 19'b1111111111111011110, 19'b1111111111111111111, 19'b1111111111111101101, 19'b0000000000000000010, 19'b0000000000000110000, 19'b0000000000000011110, 19'b0000000000001110101, 19'b0000000000000010101, 19'b1111111111111010100, 19'b0000000000000000000, 19'b0000000000000010001, 19'b1111111111111110110, 19'b0000000000001101011, 19'b0000000000001001100, 19'b0000000000000110001, 19'b1111111111111111111, 19'b1111111111110110010, 19'b1111111111111111001, 19'b0000000000000110010}, 
{19'b0000000000001000110, 19'b0000000000000001001, 19'b0000000000000011011, 19'b1111111111111111011, 19'b1111111111011111011, 19'b0000000000000000000, 19'b0000000000000000000, 19'b0000000000001110011, 19'b0000000000001111100, 19'b1111111111111111001, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000000000000, 19'b0000000000000000010, 19'b1111111111111110110, 19'b0000000000001101101, 19'b0000000000000000000, 19'b1111111111111110011, 19'b1111111111111111111, 19'b1111111111110100101, 19'b1111111111111100000, 19'b0000000000000011001, 19'b1111111111111011111, 19'b1111111111111111111, 19'b0000000000000000001, 19'b1111111111111100110, 19'b0000000000000100101, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111110010001, 19'b0000000000010011110}, 
{19'b1111111111010100010, 19'b1111111111111110011, 19'b1111111111111111101, 19'b0000000000000000010, 19'b1111111111111110010, 19'b0000000000000000011, 19'b1111111111111100110, 19'b1111111111110110011, 19'b0000000000000011011, 19'b1111111111111110101, 19'b1111111111111111001, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000001101011, 19'b0000000000000000000, 19'b0000000000010101000, 19'b1111111111111111111, 19'b0000000000001101111, 19'b1111111111100110011, 19'b0000000000000000000, 19'b1111111111111000110, 19'b0000000000001010110, 19'b0000000000010000100, 19'b0000000000000000000, 19'b0000000000000010111, 19'b0000000000001010011, 19'b0000000000001111010, 19'b0000000000000001000, 19'b1111111111111111101, 19'b1111111111111111111, 19'b1111111111111111000, 19'b0000000000001110011}, 
{19'b0000000000000011101, 19'b1111111111111111111, 19'b0000000000001001100, 19'b1111111111010110011, 19'b1111111110100111110, 19'b1111111111101001100, 19'b0000000000010110101, 19'b1111111111011000001, 19'b1111111111111111111, 19'b1111111111010100101, 19'b1111111111011111111, 19'b1111111111101010001, 19'b0000000000010110100, 19'b1111111111111111111, 19'b1111111111111111000, 19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111110111100, 19'b1111111111111111111, 19'b1111111111100000101, 19'b0000000000000000000, 19'b0000000000001011111, 19'b1111111111111111111, 19'b0000000000000001011, 19'b0000000000010001001, 19'b0000000000000011010, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000001101001, 19'b1111111111111101110, 19'b0000000000001100110}, 
{19'b1111111111111101101, 19'b1111111111110101111, 19'b1111111111110000100, 19'b1111111111111100111, 19'b1111111111101101100, 19'b0000000000000100001, 19'b1111111111110100011, 19'b1111111111110110111, 19'b1111111111100101011, 19'b0000000000000011000, 19'b1111111111111111101, 19'b1111111111110101110, 19'b0000000000000111100, 19'b1111111111111111010, 19'b1111111111111101010, 19'b1111111111011100100, 19'b1111111111111111111, 19'b0000000000000101011, 19'b0000000000001100010, 19'b1111111111110101100, 19'b1111111111110110011, 19'b1111111111111011111, 19'b1111111111111111111, 19'b0000000000000001110, 19'b1111111111111101000, 19'b1111111111010110100, 19'b1111111111101111000, 19'b1111111111111101000, 19'b0000000000000000010, 19'b1111111111111110101, 19'b0000000000000001111, 19'b1111111111111111111}, 
{19'b1111111111110110001, 19'b1111111111111010001, 19'b1111111111111010111, 19'b1111111111110000110, 19'b1111111111111000100, 19'b1111111111111111111, 19'b0000000000000110101, 19'b1111111111111010111, 19'b0000000000001100110, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111111111111, 19'b0000000000001110000, 19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111111111011011, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111111111111, 19'b0000000000000010110, 19'b1111111111110100011, 19'b0000000000000000111, 19'b1111111111111111111, 19'b1111111111111011011, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111111111111}, 
{19'b1111111111100001011, 19'b1111111111111100010, 19'b1111111111100111101, 19'b0000000000000111110, 19'b0000000000011111001, 19'b1111111111111111111, 19'b1111111111111110001, 19'b0000000000001111010, 19'b1111111111100011111, 19'b1111111111111101000, 19'b0000000000000000000, 19'b1111111111110011000, 19'b1111111111111111111, 19'b0000000000000100110, 19'b1111111111110011110, 19'b0000000000110000010, 19'b1111111111111111011, 19'b0000000000000010111, 19'b0000000000001101010, 19'b0000000000001111101, 19'b0000000000000000000, 19'b1111111111101010100, 19'b0000000000000000000, 19'b0000000000011010010, 19'b1111111111110100011, 19'b0000000000101100101, 19'b1111111111110110011, 19'b1111111111110010111, 19'b1111111111100001110, 19'b1111111111100010010, 19'b0000000000000000000, 19'b0000000000000011011}, 
{19'b0000000000000000000, 19'b1111111111111111000, 19'b1111111111111011010, 19'b0000000000000000000, 19'b0000000000010011101, 19'b1111111111111110101, 19'b1111111111111011111, 19'b0000000000000101111, 19'b0000000000000110011, 19'b0000000000000000001, 19'b1111111111111111011, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111111000101, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111111111101, 19'b0000000000000000001, 19'b0000000000000101011, 19'b0000000000000001001, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000000000011, 19'b0000000000000010011, 19'b1111111111110111100, 19'b0000000000000100010, 19'b0000000000001111111, 19'b1111111111111111111, 19'b0000000000000000011, 19'b0000000000000011001, 19'b0000000000000100011}, 
{19'b0000000000000110001, 19'b0000000000000000000, 19'b1111111111111001011, 19'b1111111111101111111, 19'b1111111111001101001, 19'b0000000000001000100, 19'b0000000000000000000, 19'b1111111111001011000, 19'b0000000000000010010, 19'b1111111111111111111, 19'b0000000000000000001, 19'b1111111111111111111, 19'b0000000000000000101, 19'b0000000000000000000, 19'b1111111111111110110, 19'b1111111111100111100, 19'b1111111111111111111, 19'b0000000000001110000, 19'b0000000000001000000, 19'b0000000000001100001, 19'b1111111111100011110, 19'b1111111111101001001, 19'b0000000000000111101, 19'b1111111111111101110, 19'b1111111111111101000, 19'b0000000000010110111, 19'b1111111111111001110, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000001101100, 19'b1111111111111111111, 19'b0000000000000000011}, 
{19'b1111111111110011010, 19'b1111111111100000011, 19'b0000000000000000000, 19'b1111111111111111110, 19'b0000000000010101010, 19'b1111111111101110110, 19'b1111111111110001110, 19'b0000000000000111011, 19'b1111111111111111111, 19'b0000000000001001100, 19'b0000000000000100101, 19'b1111111111111011001, 19'b0000000000000000000, 19'b0000000000000000111, 19'b1111111111111110101, 19'b1111111111101111110, 19'b0000000000001011001, 19'b0000000000000001110, 19'b0000000000010011000, 19'b0000000000000101100, 19'b0000000000000000000, 19'b1111111111111101100, 19'b0000000000001000000, 19'b1111111111111010011, 19'b1111111111101100010, 19'b1111111111111111100, 19'b0000000000001011110, 19'b1111111111111111111, 19'b0000000000000000100, 19'b1111111111111001111, 19'b0000000000001000110, 19'b0000000000010001101}, 
{19'b0000000000000000111, 19'b0000000000000000000, 19'b0000000000001110000, 19'b0000000000000000100, 19'b1111111111111101011, 19'b0000000000001011100, 19'b0000000000000101111, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111110111000, 19'b1111111111111100100, 19'b1111111111110101010, 19'b1111111111111111111, 19'b0000000000000011001, 19'b1111111111111011100, 19'b0000000000110101111, 19'b0000000000000000000, 19'b1111111111111001111, 19'b1111111111110011111, 19'b1111111111111111001, 19'b0000000000001100101, 19'b0000000000001000001, 19'b0000000000000000000, 19'b1111111111111111110, 19'b0000000000001110000, 19'b0000000000010001001, 19'b0000000000011111101, 19'b0000000000000000101, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111111111001, 19'b1111111111111011011}, 
{19'b1111111111110110000, 19'b0000000000000011000, 19'b0000000000000010100, 19'b1111111111110000001, 19'b1111111111101110110, 19'b0000000000011110000, 19'b0000000000000011001, 19'b0000000000000000000, 19'b1111111111110101101, 19'b1111111111111010010, 19'b0000000000001000010, 19'b0000000000000100100, 19'b0000000000000000000, 19'b1111111111111010111, 19'b0000000000010010010, 19'b1111111111111111111, 19'b1111111111111111001, 19'b0000000000000000000, 19'b0000000000000000110, 19'b1111111111111101000, 19'b0000000000000101000, 19'b0000000000000001000, 19'b0000000000000111010, 19'b1111111111111111111, 19'b0000000000000000001, 19'b0000000000101010000, 19'b1111111111111100011, 19'b1111111111111110100, 19'b1111111111111111111, 19'b1111111111111001000, 19'b1111111111111101011, 19'b0000000000001011010}, 
{19'b0000000000000011110, 19'b0000000000000100101, 19'b0000000000010100111, 19'b1111111111111101011, 19'b0000000000000110011, 19'b0000000000010110011, 19'b0000000000000000000, 19'b1111111111111110000, 19'b0000000000000111100, 19'b1111111111111000101, 19'b1111111111111111111, 19'b1111111111111000010, 19'b0000000000000000000, 19'b0000000000011001001, 19'b1111111111111110110, 19'b0000000000000000000, 19'b0000000000001111000, 19'b0000000000000000000, 19'b0000000000000000001, 19'b1111111111101011111, 19'b1111111111110000010, 19'b1111111111111101101, 19'b1111111111111111111, 19'b1111111111110110101, 19'b1111111111111101101, 19'b1111111111111010101, 19'b1111111111110011011, 19'b1111111111110010011, 19'b0000000000000001111, 19'b0000000000000111001, 19'b1111111111100110100, 19'b0000000000000000001}, 
{19'b1111111111101100111, 19'b0000000000000000000, 19'b1111111111111111000, 19'b1111111111111100110, 19'b1111111111111111111, 19'b0000000000001000100, 19'b1111111111111011000, 19'b0000000000010001010, 19'b1111111111101000110, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111111111110, 19'b1111111111111010001, 19'b0000000000000101000, 19'b0000000000001011101, 19'b1111111111111111011, 19'b1111111111101111111, 19'b1111111111111100001, 19'b0000000000000111001, 19'b0000000000000100000, 19'b0000000000000000000, 19'b0000000000000000001, 19'b0000000000000101001, 19'b1111111111110000101, 19'b0000000000000000000, 19'b1111111111111111111, 19'b0000000000000000001, 19'b0000000000000000000, 19'b1111111111110111111}, 
{19'b1111111111101010011, 19'b1111111111111111101, 19'b1111111111111111110, 19'b1111111111111110111, 19'b1111111111111111101, 19'b0000000000000110110, 19'b0000000000000000011, 19'b0000000000000010001, 19'b0000000000000010011, 19'b0000000000000100000, 19'b0000000000000101000, 19'b0000000000001010010, 19'b0000000000000001101, 19'b1111111111111001110, 19'b0000000000000000000, 19'b0000000000011000011, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111111111110, 19'b0000000000000111000, 19'b0000000000001001000, 19'b0000000000000001111, 19'b0000000000000010101, 19'b1111111111111110000, 19'b1111111111111101111, 19'b0000000000000001101, 19'b1111111111111011101, 19'b1111111111110111111, 19'b0000000000001101011, 19'b1111111111111110000, 19'b0000000000000010000, 19'b1111111111110011111}, 
{19'b0000000000000000000, 19'b1111111111111111111, 19'b0000000000000010011, 19'b0000000000000000000, 19'b0000000000111010000, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111111111111, 19'b0000000000000111000, 19'b1111111111111011001, 19'b0000000000000000000, 19'b0000000000000000000, 19'b0000000000000000000, 19'b0000000000001000010, 19'b0000000000000000000, 19'b1111111111110110101, 19'b1111111111111111111, 19'b1111111111111011101, 19'b0000000000010100111, 19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000000100010, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000000010101}, 
{19'b1111111111111111110, 19'b0000000000000001110, 19'b1111111111111111111, 19'b0000000000000011000, 19'b1111111111111101001, 19'b1111111111111000010, 19'b1111111111111100000, 19'b0000000000010001110, 19'b0000000000000000000, 19'b0000000000000110001, 19'b1111111111111111010, 19'b0000000000000100001, 19'b1111111111111101111, 19'b1111111111110101111, 19'b1111111111110011110, 19'b0000000000000000110, 19'b1111111111111111111, 19'b1111111111111101110, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111111111111, 19'b0000000000000100110, 19'b0000000000000010010, 19'b1111111111110111111, 19'b0000000000000111001, 19'b1111111111110101011, 19'b0000000000000000001, 19'b0000000000000000000, 19'b1111111111110101010, 19'b0000000000000000000, 19'b0000000000000010111, 19'b1111111111111110000}, 
{19'b1111111111111111010, 19'b1111111111111001101, 19'b0000000000000000000, 19'b1111111111111100001, 19'b0000000000001101110, 19'b1111111111111111111, 19'b1111111111111110101, 19'b0000000000000110110, 19'b1111111111100110111, 19'b0000000000000000000, 19'b1111111111111101100, 19'b1111111111111111110, 19'b0000000000010110011, 19'b0000000000001110101, 19'b1111111111111001101, 19'b1111111111111110101, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111110111010, 19'b1111111111111000011, 19'b0000000000001000011, 19'b0000000000000000000, 19'b1111111111110111001, 19'b0000000000000001100, 19'b1111111111111010110, 19'b1111111111111101110, 19'b0000000000001000101, 19'b0000000000000000000, 19'b1111111111110000001}, 
{19'b0000000000101000100, 19'b0000000000010101111, 19'b1111111111110000000, 19'b0000000000000000001, 19'b1111111111101001110, 19'b0000000000000000000, 19'b0000000000001110010, 19'b0000000000000001111, 19'b0000000000001110010, 19'b1111111111111111111, 19'b1111111111110110000, 19'b1111111111111010111, 19'b0000000000001001000, 19'b0000000000000001110, 19'b1111111111111001101, 19'b0000000000001000011, 19'b0000000000100010010, 19'b1111111111110111101, 19'b1111111111101101000, 19'b0000000000000000000, 19'b1111111111111110001, 19'b1111111111110100101, 19'b1111111111111111001, 19'b1111111111111111111, 19'b0000000000000101100, 19'b1111111111101000111, 19'b0000000000000101101, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000000110111, 19'b1111111111111110001, 19'b0000000000000011110}, 
{19'b1111111111111010000, 19'b1111111111110011101, 19'b1111111111111101101, 19'b1111111111110101010, 19'b1111111111111110111, 19'b0000000000000011001, 19'b0000000000000000000, 19'b1111111111111111010, 19'b0000000000000010011, 19'b1111111111111111110, 19'b0000000000000000000, 19'b1111111111110010000, 19'b0000000000000110100, 19'b0000000000000101001, 19'b1111111111111001011, 19'b0000000000011100011, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111111111101, 19'b0000000000000000000, 19'b0000000000010100001, 19'b1111111111100001111, 19'b1111111111111001000, 19'b1111111111111100011, 19'b1111111111111110110, 19'b0000000000001100100, 19'b1111111111111100101, 19'b0000000000000001001, 19'b0000000000011110111, 19'b1111111111011111001, 19'b1111111111101000100, 19'b0000000000000001011}, 
{19'b0000000000000001000, 19'b1111111111111100001, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111010001111, 19'b1111111111011001001, 19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111111101111000, 19'b0000000000000001100, 19'b0000000000000000000, 19'b1111111111111110001, 19'b0000000000000000000, 19'b1111111111111100010, 19'b1111111111111100101, 19'b1111111111111011100, 19'b1111111111110110100, 19'b0000000000010010000, 19'b0000000000000000000, 19'b0000000000000010111, 19'b1111111111111111111, 19'b1111111111111011011, 19'b0000000000000000000, 19'b1111111111111010011, 19'b0000000000001110000, 19'b1111111111011000001, 19'b0000000000001110000, 19'b1111111111111111111, 19'b1111111111111111101, 19'b0000000000001100110, 19'b1111111111111111111, 19'b0000000000001111000}, 
{19'b1111111111111111111, 19'b0000000000000000010, 19'b1111111111111101001, 19'b0000000000000100110, 19'b0000000000000011100, 19'b1111111111101010000, 19'b0000000000000000000, 19'b0000000000000100000, 19'b0000000000100101000, 19'b1111111111111111011, 19'b0000000000000000000, 19'b0000000000000011100, 19'b0000000000010110111, 19'b1111111111111101111, 19'b0000000000000000111, 19'b0000000000000110011, 19'b1111111111111111111, 19'b0000000000000001110, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111101110011, 19'b0000000000000010011, 19'b0000000000000100011, 19'b0000000000000001011, 19'b1111111111111111111, 19'b0000000000001101111, 19'b0000000000000000010, 19'b0000000000001000000, 19'b1111111111100101010, 19'b0000000000000110100, 19'b0000000000011001010, 19'b0000000000000000010}, 
{19'b1111111111101001100, 19'b0000000000001101100, 19'b1111111111101111010, 19'b0000000000000111110, 19'b1111111111111001010, 19'b0000000000000000000, 19'b0000000000011111110, 19'b1111111111110001000, 19'b1111111111101101010, 19'b0000000000001010111, 19'b1111111111110001101, 19'b1111111111111110011, 19'b1111111111111111111, 19'b0000000000010110000, 19'b1111111111111111111, 19'b1111111111101100101, 19'b1111111111111111111, 19'b0000000000011100001, 19'b1111111111100001110, 19'b1111111111111110011, 19'b0000000000010100010, 19'b1111111111101000110, 19'b0000000000000011011, 19'b1111111111111111000, 19'b0000000000010001010, 19'b1111111111011111011, 19'b1111111111101000110, 19'b1111111111110011011, 19'b1111111111111111111, 19'b0000000000000110101, 19'b0000000000000001100, 19'b0000000000001011011}, 
{19'b1111111111111010001, 19'b0000000000000011010, 19'b1111111111111111111, 19'b0000000000001001100, 19'b1111111111111101100, 19'b0000000000001110100, 19'b0000000000000000001, 19'b1111111111111111010, 19'b1111111111111111110, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000100001010, 19'b0000000000000000110, 19'b0000000000001100000, 19'b0000000000000000000, 19'b1111111111110010011, 19'b1111111111111011000, 19'b1111111111111111111, 19'b1111111111111110111, 19'b0000000000000010101, 19'b1111111111111111111, 19'b1111111111110100001, 19'b1111111111111111111, 19'b0000000000010010111, 19'b0000000000010011110, 19'b1111111111111111111, 19'b1111111111111110111, 19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111111111001110}, 
{19'b1111111111111010110, 19'b0000000000000000000, 19'b0000000000010001011, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111111000101, 19'b0000000000000000000, 19'b1111111111001000101, 19'b0000000000001101110, 19'b0000000000000000111, 19'b0000000000000001101, 19'b1111111111101000111, 19'b0000000000000000001, 19'b1111111111110111001, 19'b1111111111111101111, 19'b0000000000000000000, 19'b0000000000000001010, 19'b0000000000000000000, 19'b0000000000000111001, 19'b0000000000000000000, 19'b1111111111111111011, 19'b0000000000010101000, 19'b0000000000011000000, 19'b1111111111110001110, 19'b1111111111110110111, 19'b0000000000001111111, 19'b1111111111101100011, 19'b0000000000000001111, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000001011110}, 
{19'b1111111111111000101, 19'b1111111111111111111, 19'b1111111111110000101, 19'b1111111111110011000, 19'b1111111111111111000, 19'b1111111111110111010, 19'b0000000000000000000, 19'b0000000000000101110, 19'b1111111111110000101, 19'b1111111111111010101, 19'b1111111111111100110, 19'b0000000000000000000, 19'b0000000000000001110, 19'b1111111111111111010, 19'b1111111111111100000, 19'b0000000000000110000, 19'b0000000000001110010, 19'b0000000000001000011, 19'b1111111111110111101, 19'b0000000000000011000, 19'b1111111111111111001, 19'b1111111111111110001, 19'b0000000000000001011, 19'b0000000000000001000, 19'b1111111111111011100, 19'b0000000000000101101, 19'b1111111111111010001, 19'b0000000000000011110, 19'b1111111111111111111, 19'b1111111111101101000, 19'b1111111111111110010, 19'b0000000000001110011}, 
{19'b1111111111111110010, 19'b1111111111111010101, 19'b0000000000000100111, 19'b0000000000010000001, 19'b0000000000000101011, 19'b0000000000000101010, 19'b0000000000000010111, 19'b1111111111110011000, 19'b1111111111110010110, 19'b0000000000000100011, 19'b0000000000000000110, 19'b0000000000000010110, 19'b0000000000000001011, 19'b0000000000000000010, 19'b0000000000001101001, 19'b0000000000000000011, 19'b1111111111111100100, 19'b0000000000000110100, 19'b1111111111111110000, 19'b1111111111111101101, 19'b0000000000000111000, 19'b1111111111111000000, 19'b1111111111111110010, 19'b0000000000001000001, 19'b0000000000000001011, 19'b1111111111111001001, 19'b1111111111110011010, 19'b1111111111111111001, 19'b1111111111101110001, 19'b0000000000000011110, 19'b0000000000000110100, 19'b0000000000000000000}, 
{19'b1111111111111111001, 19'b1111111111111110101, 19'b1111111111111111001, 19'b1111111111111101110, 19'b1111111111110111100, 19'b1111111111110111000, 19'b0000000000000100000, 19'b0000000000000000100, 19'b1111111111110100010, 19'b0000000000001010101, 19'b1111111111111110101, 19'b1111111111111111111, 19'b1111111111111000111, 19'b0000000000000000010, 19'b0000000000000001111, 19'b1111111111111100101, 19'b1111111111111110111, 19'b1111111111111101010, 19'b1111111111111010110, 19'b0000000000000000000, 19'b1111111111110111000, 19'b0000000000000110100, 19'b1111111111110010011, 19'b0000000000000000010, 19'b0000000000000010101, 19'b0000000000000111111, 19'b0000000000000001101, 19'b0000000000000000011, 19'b0000000000010010101, 19'b0000000000000011010, 19'b0000000000000000000, 19'b0000000000000101010}, 
{19'b1111111111111110110, 19'b0000000000010000001, 19'b1111111111111111111, 19'b1111111111111101111, 19'b1111111111110010010, 19'b1111111111111011001, 19'b0000000000011010010, 19'b1111111111010011111, 19'b1111111111101001101, 19'b1111111111110011001, 19'b1111111111110001111, 19'b1111111111101111110, 19'b1111111111111111111, 19'b0000000000011110111, 19'b1111111111111110010, 19'b0000000000000000000, 19'b1111111111110010011, 19'b0000000000011100100, 19'b1111111111100101100, 19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111111101010011, 19'b0000000000000000000, 19'b1111111111111111111, 19'b0000000000000011100, 19'b1111111111111100010, 19'b1111111111110110100, 19'b1111111111111111111, 19'b0000000000001011001, 19'b0000000000000000001, 19'b1111111111111010110, 19'b0000000000000000000}, 
{19'b0000000000010111100, 19'b1111111111111000110, 19'b0000000000001000011, 19'b1111111111111101111, 19'b0000000000000100111, 19'b1111111111111111110, 19'b1111111111111111110, 19'b1111111111111010000, 19'b0000000000000000000, 19'b0000000000000101111, 19'b1111111111111111111, 19'b1111111111111100001, 19'b1111111111111111111, 19'b0000000000001110101, 19'b0000000000000001001, 19'b0000000000000010100, 19'b0000000000000001100, 19'b1111111111111110011, 19'b0000000000000001010, 19'b0000000000000000000, 19'b1111111111111111011, 19'b1111111111111111111, 19'b1111111111101100011, 19'b1111111111111111111, 19'b0000000000000011101, 19'b1111111111111000100, 19'b1111111111110111010, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000100011101, 19'b1111111111101101101, 19'b1111111111111000100}, 
{19'b1111111111111101001, 19'b1111111111111001011, 19'b1111111111111011110, 19'b0000000000000010010, 19'b0000000000001000111, 19'b1111111111110111101, 19'b1111111111111111111, 19'b1111111111110001111, 19'b0000000000000011111, 19'b0000000000001000101, 19'b1111111111110010010, 19'b1111111111101111110, 19'b0000000000000001100, 19'b1111111111010100010, 19'b1111111111111011001, 19'b1111111111111000000, 19'b1111111111110011010, 19'b1111111111111111111, 19'b0000000000001000100, 19'b0000000000000000000, 19'b1111111111111101000, 19'b1111111111111101001, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111111100001, 19'b1111111111001111101, 19'b1111111111011100011, 19'b1111111111101110100, 19'b0000000000000011100, 19'b0000000000001101001, 19'b1111111111111111111, 19'b0000000000001111011}, 
{19'b1111111111111010000, 19'b1111111111110010010, 19'b0000000000001010011, 19'b0000000000000100110, 19'b0000000000000010110, 19'b1111111111111010000, 19'b1111111111111101111, 19'b0000000000000110010, 19'b0000000000100010011, 19'b1111111111110101000, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000000111100, 19'b1111111111111100011, 19'b1111111111111110110, 19'b1111111111111110111, 19'b1111111111111001100, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000001110100, 19'b1111111111110111011, 19'b1111111111111111110, 19'b0000000000001000001, 19'b1111111111111111010, 19'b0000000000000000000, 19'b0000000000100001101, 19'b0000000000010100110, 19'b0000000000000000001, 19'b0000000000000000000, 19'b1111111111100101000, 19'b1111111111111011101, 19'b1111111111111111111}, 
{19'b0000000000000000111, 19'b0000000000000011000, 19'b1111111111111111000, 19'b0000000000000000000, 19'b0000000000001110110, 19'b1111111111100001000, 19'b0000000000000000000, 19'b1111111111111001111, 19'b0000000000001011111, 19'b0000000000000000000, 19'b1111111111111110110, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111111111111, 19'b0000000000000000010, 19'b1111111111111001000, 19'b0000000000010000100, 19'b1111111111111111101, 19'b1111111111111111000, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111111111100, 19'b0000000000000000000, 19'b1111111111111111111, 19'b0000000000000000110, 19'b1111111111101011101, 19'b0000000000000011010, 19'b0000000000001011101, 19'b1111111111111111110, 19'b0000000000000110000, 19'b1111111111111111111, 19'b0000000000000100110}, 
{19'b1111111111110011000, 19'b0000000000000000100, 19'b1111111111100001001, 19'b0000000000000000011, 19'b1111111111111100110, 19'b1111111111111101011, 19'b1111111111111111111, 19'b1111111111111010001, 19'b1111111111111101101, 19'b1111111111111011110, 19'b0000000000000011000, 19'b0000000000000001101, 19'b1111111111110100101, 19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111111111111011, 19'b0000000000000100100, 19'b1111111111111110101, 19'b1111111111111110001, 19'b1111111111111110001, 19'b1111111111111111111, 19'b0000000000010001010, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111111111011, 19'b0000000000010100010, 19'b0000000000001100000, 19'b0000000000000010001, 19'b1111111111111001110, 19'b1111111111111111010, 19'b0000000000000100001, 19'b0000000000000011101}, 
{19'b0000000000000010001, 19'b0000000000000010100, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111100010000, 19'b0000000000000010110, 19'b0000000000000001100, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111110101001, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111110101101, 19'b0000000000000000000, 19'b0000000000000000000, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111101001001, 19'b0000000000000000100, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000001000010, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000011101001, 19'b0000000000010101110, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111110001000, 19'b0000000000000000000, 19'b1111111111111111111}, 
{19'b0000000000000100110, 19'b0000000000000011011, 19'b0000000000010000001, 19'b1111111111110000000, 19'b0000000000001000011, 19'b0000000000000111100, 19'b0000000000000000011, 19'b0000000000001100010, 19'b0000000000000000110, 19'b1111111111111111001, 19'b0000000000000010011, 19'b0000000000000000010, 19'b1111111111111111111, 19'b0000000000000111101, 19'b1111111111111111101, 19'b1111111111111101011, 19'b0000000000000000000, 19'b0000000000000010000, 19'b1111111111111100111, 19'b0000000000000110010, 19'b0000000000000010000, 19'b1111111111011010110, 19'b1111111111111000101, 19'b0000000000000101110, 19'b1111111111111111111, 19'b1111111111011111101, 19'b1111111111110111111, 19'b1111111111111110100, 19'b1111111111111111111, 19'b1111111111111100010, 19'b0000000000000000000, 19'b1111111111111101011}, 
{19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111111111010001, 19'b1111111111110101001, 19'b0000000000000010101, 19'b0000000000000000000, 19'b0000000000000110000, 19'b1111111111111111101, 19'b0000000000001111111, 19'b1111111111111111101, 19'b0000000000000000000, 19'b1111111111101010000, 19'b1111111111111111111, 19'b0000000000001000000, 19'b1111111111111111111, 19'b1111111111101111010, 19'b0000000000000000000, 19'b1111111111111111010, 19'b0000000000010000110, 19'b1111111111111111111, 19'b1111111111100100000, 19'b1111111111111111111, 19'b0000000000010000100, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000001000111, 19'b1111111111111001111, 19'b0000000000000100011, 19'b0000000000000000000, 19'b1111111111110011000, 19'b0000000000000000000, 19'b0000000000000000001}, 
{19'b1111111111110010001, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111111111100, 19'b0000000000011111101, 19'b1111111111111000000, 19'b1111111111111111101, 19'b1111111111111111100, 19'b1111111111111101001, 19'b1111111111111100110, 19'b0000000000000100001, 19'b0000000000001000100, 19'b1111111111111101101, 19'b0000000000001111111, 19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111111101101110, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111111010111, 19'b0000000000000000001, 19'b0000000000000010011, 19'b0000000000000000110, 19'b1111111111111111011, 19'b1111111111111100101, 19'b1111111111110011000, 19'b1111111111101101000, 19'b0000000000000000000, 19'b1111111111111000110, 19'b0000000000000010100, 19'b1111111111111111111, 19'b0000000000000100110}, 
{19'b1111111111100101100, 19'b1111111111110101111, 19'b1111111111110110000, 19'b0000000000000000000, 19'b0000000000100100100, 19'b1111111111110001110, 19'b0000000000000000000, 19'b1111111111111100100, 19'b1111111111100101110, 19'b0000000000001000110, 19'b1111111111111111111, 19'b0000000000100100010, 19'b0000000000000000000, 19'b1111111111111100111, 19'b1111111111111111111, 19'b0000000000000010000, 19'b1111111111111110110, 19'b0000000000000000000, 19'b1111111111111101000, 19'b0000000000011111101, 19'b0000000000000010011, 19'b1111111111111101010, 19'b0000000000000111000, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111111001110, 19'b1111111111111101000, 19'b1111111111100010000, 19'b1111111111110110110, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111111100001}, 
{19'b0000000000001110011, 19'b1111111111001100110, 19'b1111111111010001101, 19'b1111111111110101000, 19'b0000000000101010110, 19'b1111111111111111111, 19'b1111111111101001110, 19'b0000000000010000111, 19'b0000000000000011110, 19'b0000000000000000000, 19'b0000000000001101010, 19'b1111111111101110101, 19'b0000000000000000000, 19'b0000000000000000010, 19'b1111111111111101111, 19'b0000000000000001001, 19'b1111111111111001010, 19'b1111111111000101000, 19'b0000000000001010101, 19'b0000000000010110000, 19'b0000000000010000111, 19'b0000000000000000001, 19'b0000000000000001110, 19'b1111111111100110001, 19'b1111111111010111100, 19'b1111111111111111101, 19'b1111111111101100110, 19'b1111111111100010101, 19'b1111111111110011100, 19'b1111111111000111110, 19'b0000000000011010110, 19'b0000000000011011011}, 
{19'b0000000000000000000, 19'b0000000000000000000, 19'b0000000000000000001, 19'b0000000000000000000, 19'b0000000000010000100, 19'b1111111111110100000, 19'b0000000000000001001, 19'b0000000000000100101, 19'b1111111111101001101, 19'b0000000000000010010, 19'b1111111111111111101, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000001111010, 19'b0000000000000011010, 19'b0000000000000001011, 19'b0000000000000011111, 19'b0000000000010101010, 19'b1111111111110010000, 19'b0000000000000000000, 19'b1111111111110101011, 19'b1111111111111111111, 19'b0000000000010100001, 19'b0000000000000000100, 19'b1111111111111111110, 19'b1111111111011100000, 19'b1111111111111111011, 19'b1111111111110110000, 19'b1111111111111100000, 19'b0000000000000000001, 19'b0000000000001000101, 19'b0000000000000110101}, 
{19'b1111111111111101001, 19'b0000000000001000100, 19'b1111111111101100100, 19'b0000000000000001010, 19'b0000000000001100011, 19'b1111111111111101011, 19'b1111111111111111101, 19'b0000000000001010011, 19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111111111011110, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111111101110, 19'b1111111111111000001, 19'b1111111111111011110, 19'b1111111111111100011, 19'b1111111111111011111, 19'b1111111111111000111, 19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111111111101001, 19'b1111111111111011101, 19'b0000000000011001011, 19'b0000000000000000000, 19'b1111111111101000111, 19'b1111111111111111011, 19'b0000000000000111111, 19'b0000000000000000000, 19'b0000000000000000000, 19'b0000000000010000000, 19'b1111111111111111111}, 
{19'b1111111111111111111, 19'b0000000000000000010, 19'b1111111111111111111, 19'b1111111111110110000, 19'b1111111111001000111, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111111111100, 19'b1111111111011001101, 19'b0000000000000101001, 19'b1111111111111001101, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111101000010, 19'b1111111111111101000, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000000000100, 19'b0000000000000010010, 19'b0000000000010110000, 19'b1111111111111000010, 19'b1111111111101100110, 19'b0000000000000000000, 19'b1111111111101111011, 19'b1111111111111001101, 19'b1111111111110001001, 19'b1111111111111111100, 19'b1111111111111111001, 19'b1111111111111110110, 19'b1111111111100001110, 19'b1111111111111101110, 19'b0000000000001111100}, 
{19'b0000000000000111001, 19'b0000000000001110000, 19'b1111111111111111110, 19'b0000000000001010001, 19'b1111111111110010100, 19'b1111111111111000000, 19'b0000000000000110000, 19'b0000000000000100011, 19'b1111111111111100111, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111101011011, 19'b1111111111111111111, 19'b0000000000001001001, 19'b1111111111111000101, 19'b0000000000000010001, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000001101010, 19'b1111111111101011000, 19'b0000000000010001111, 19'b0000000000000011000, 19'b0000000000000000000, 19'b0000000000001101100, 19'b0000000000000000001, 19'b1111111111111101101, 19'b1111111111100111101, 19'b1111111111111000111, 19'b1111111111110101000, 19'b0000000000001011010}, 
{19'b0000000000000000000, 19'b0000000000000000011, 19'b1111111111101000100, 19'b1111111111111111110, 19'b0000000000001101001, 19'b1111111111110110111, 19'b1111111111111111001, 19'b1111111111111111111, 19'b0000000000000001010, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111110010111, 19'b0000000000000110001, 19'b0000000000000000011, 19'b0000000000000000000, 19'b0000000000000010011, 19'b1111111111111111111, 19'b1111111111110110011, 19'b0000000000000001001, 19'b0000000000000000000, 19'b1111111111111101110, 19'b1111111111111110100, 19'b0000000000010010111, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111101101010, 19'b1111111111101011000, 19'b0000000000001111011, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000000001110, 19'b0000000000010010000}, 
{19'b1111111111101010001, 19'b1111111111111111111, 19'b1111111111110010011, 19'b0000000000000000010, 19'b1111111111101001011, 19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111111111011110, 19'b1111111111011101111, 19'b1111111111111110010, 19'b0000000000000000000, 19'b1111111111111111011, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111111111011, 19'b1111111111111100110, 19'b1111111111110110100, 19'b1111111111111001111, 19'b0000000000000100001, 19'b1111111111111111110, 19'b1111111111111110011, 19'b0000000000000000000, 19'b0000000000010101100, 19'b1111111111111111111, 19'b0000000000001001100, 19'b0000000000000101110, 19'b1111111111110111001, 19'b0000000000001101101, 19'b1111111111111101000, 19'b0000000000000000000, 19'b1111111111111111111, 19'b0000000000100101010}, 
{19'b1111111111101011111, 19'b0000000000000001111, 19'b0000000000000011001, 19'b1111111111111110001, 19'b0000000000001111101, 19'b1111111111101100101, 19'b1111111111111111100, 19'b0000000000010000111, 19'b0000000000001010001, 19'b0000000000000000100, 19'b1111111111111111111, 19'b1111111111111011100, 19'b1111111111111010010, 19'b1111111111111011110, 19'b1111111111111100110, 19'b0000000000000101110, 19'b1111111111111111111, 19'b0000000000000000100, 19'b0000000000001001000, 19'b0000000000000000000, 19'b0000000000000000000, 19'b0000000000000000111, 19'b0000000000010000001, 19'b0000000000000010111, 19'b0000000000000000011, 19'b1111111111111001000, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111111111000, 19'b1111111111111111001, 19'b1111111111111111111, 19'b0000000000000100010}, 
{19'b1111111111111111111, 19'b0000000000000000001, 19'b1111111111110010011, 19'b1111111111111011001, 19'b0000000000010010000, 19'b1111111111111111111, 19'b1111111111111011000, 19'b0000000000001111101, 19'b1111111111111100100, 19'b0000000000010010101, 19'b0000000000000101011, 19'b1111111111111000010, 19'b0000000000000000000, 19'b0000000000000000001, 19'b1111111111111111000, 19'b0000000000000001010, 19'b1111111111111011000, 19'b1111111111101111001, 19'b0000000000010001110, 19'b0000000000001001111, 19'b0000000000101000100, 19'b0000000000001100110, 19'b0000000000001111111, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000000000000, 19'b0000000000000011101, 19'b0000000000000101000, 19'b1111111111100101000, 19'b1111111111111111111, 19'b1111111111111111101, 19'b1111111111111111100}, 
{19'b0000000000000000000, 19'b1111111111111010011, 19'b1111111111111001010, 19'b0000000000000000000, 19'b1111111111110000011, 19'b0000000000000000000, 19'b0000000000001100010, 19'b0000000000000110111, 19'b0000000000000011011, 19'b1111111111111001101, 19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111111101010, 19'b0000000000001100111, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111101100101, 19'b0000000000000000000, 19'b1111111111110011101, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111111111101, 19'b0000000000000000111, 19'b0000000000000001000, 19'b0000000000000001110, 19'b0000000000001000110, 19'b1111111111111011110, 19'b1111111111111111100, 19'b1111111111100011010, 19'b0000000000000101000}, 
{19'b0000000000011100010, 19'b1111111111111111011, 19'b0000000000000100001, 19'b1111111111111001010, 19'b1111111111111010100, 19'b0000000000000010001, 19'b0000000000001010010, 19'b0000000000000000000, 19'b0000000000100001101, 19'b0000000000000000000, 19'b1111111111111110101, 19'b0000000000000001001, 19'b0000000000000110000, 19'b1111111111111111110, 19'b0000000000000011011, 19'b0000000000000110100, 19'b1111111111111111101, 19'b1111111111100011100, 19'b1111111111111100011, 19'b1111111111111111111, 19'b0000000000000111011, 19'b0000000000000000000, 19'b1111111111111111111, 19'b0000000000000111001, 19'b0000000000000001001, 19'b1111111111101111001, 19'b1111111111111001011, 19'b0000000000001000011, 19'b1111111111111110001, 19'b0000000000010000100, 19'b1111111111111111111, 19'b1111111111110100100}, 
{19'b0000000000000000110, 19'b0000000000000110100, 19'b1111111111111111111, 19'b1111111111111101100, 19'b1111111111101001011, 19'b1111111111111111111, 19'b0000000000000010111, 19'b1111111111111101000, 19'b0000000000001010100, 19'b1111111111111101110, 19'b1111111111111111111, 19'b1111111111111101110, 19'b1111111111111111111, 19'b1111111111111101101, 19'b0000000000000000000, 19'b0000000000010100000, 19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000000010001, 19'b0000000000001000000, 19'b0000000000000000000, 19'b0000000000000000010, 19'b0000000000000010000, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000000001010, 19'b0000000000000000000, 19'b0000000000000110001}, 
{19'b1111111111101100001, 19'b0000000000001000010, 19'b0000000000000001001, 19'b1111111111111001010, 19'b1111111111100110011, 19'b1111111111111110110, 19'b0000000000000100010, 19'b1111111111100110100, 19'b0000000000100000101, 19'b0000000000000100100, 19'b0000000000000001000, 19'b0000000000000110000, 19'b0000000000000010110, 19'b0000000000000000000, 19'b0000000000011010000, 19'b1111111111111010100, 19'b0000000000000000010, 19'b0000000000000000000, 19'b1111111111111111100, 19'b0000000000000000001, 19'b1111111111100100010, 19'b0000000000000001000, 19'b0000000000001001110, 19'b0000000000000010011, 19'b0000000000000010010, 19'b1111111111010101111, 19'b1111111111101010001, 19'b1111111111110000100, 19'b0000000000000000001, 19'b1111111111111111111, 19'b0000000000010100110, 19'b1111111111110010111}, 
{19'b1111111111111111001, 19'b1111111111110011100, 19'b1111111111111001011, 19'b1111111111100101110, 19'b1111111111101111010, 19'b0000000000010101100, 19'b0000000000010011110, 19'b1111111111110101000, 19'b0000000000000010101, 19'b1111111111111101100, 19'b1111111111111001111, 19'b1111111111101111111, 19'b0000000000000110100, 19'b1111111111101101110, 19'b0000000000001100000, 19'b1111111111111111111, 19'b0000000000010101011, 19'b1111111111111111111, 19'b1111111111111111100, 19'b1111111111110111010, 19'b1111111111111101010, 19'b1111111111111011110, 19'b1111111111101110111, 19'b0000000000000101010, 19'b1111111111111111111, 19'b1111111111111111100, 19'b1111111111110001011, 19'b0000000000010100001, 19'b0000000000010001110, 19'b1111111111111010001, 19'b1111111111010111101, 19'b0000000000001001001}, 
{19'b0000000000000000000, 19'b1111111111111110010, 19'b1111111111111111111, 19'b1111111111111001110, 19'b0000000000000001110, 19'b0000000000000000100, 19'b0000000000000100011, 19'b0000000000000000010, 19'b0000000000000111100, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000000110000, 19'b0000000000000000000, 19'b0000000000000000110, 19'b1111111111110111100, 19'b1111111111111001000, 19'b0000000000000000000, 19'b0000000000001011101, 19'b0000000000000011101, 19'b0000000000001000000, 19'b1111111111111110111, 19'b1111111111110101110, 19'b1111111111111111111, 19'b0000000000000100110, 19'b1111111111111111111, 19'b0000000000000010000, 19'b1111111111111111101, 19'b0000000000000100010, 19'b0000000000000000000, 19'b0000000000000101010, 19'b1111111111100111101, 19'b1111111111111111111}, 
{19'b0000000000010011110, 19'b1111111111111111011, 19'b0000000000001001100, 19'b1111111111101100011, 19'b1111111111110011101, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000000001110, 19'b0000000000000000001, 19'b1111111111110111111, 19'b0000000000000000000, 19'b0000000000000000001, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111110111101, 19'b0000000000001001001, 19'b1111111111111111111, 19'b1111111111111110000, 19'b0000000000000000000, 19'b0000000000000111101, 19'b1111111111110011001, 19'b0000000000000111011, 19'b0000000000001000111, 19'b0000000000001000010, 19'b1111111111111111111, 19'b0000000000100011010, 19'b1111111111110110001, 19'b0000000000010111010, 19'b1111111111111100101, 19'b1111111111101000111, 19'b1111111111110100111, 19'b0000000000001000111}, 
{19'b1111111111011101001, 19'b1111111111111110010, 19'b1111111111110110001, 19'b1111111111111111111, 19'b0000000000010000101, 19'b1111111111110100100, 19'b1111111111111100001, 19'b0000000000001111001, 19'b0000000000000110000, 19'b1111111111110000110, 19'b0000000000000000000, 19'b1111111111111110001, 19'b1111111111111111010, 19'b0000000000001000110, 19'b1111111111110000010, 19'b1111111111111111010, 19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111111111110111, 19'b0000000000000000000, 19'b1111111111110011110, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111101010111, 19'b0000000000000100011, 19'b0000000000100111101, 19'b0000000000010110001, 19'b1111111111111101101, 19'b1111111111110101101, 19'b1111111111100011010, 19'b0000000000000000000, 19'b1111111111111100111}, 
{19'b0000000000000001010, 19'b0000000000001101101, 19'b0000000000000001010, 19'b1111111111110110010, 19'b0000000000000000010, 19'b1111111111111110010, 19'b0000000000000000000, 19'b0000000000001101010, 19'b0000000000001101110, 19'b1111111111110111011, 19'b0000000000001000111, 19'b0000000000000001100, 19'b1111111111111111111, 19'b1111111111111111000, 19'b1111111111110101110, 19'b0000000000010000001, 19'b1111111111111101010, 19'b1111111111101011010, 19'b0000000000000111010, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000000111011, 19'b1111111111111011001, 19'b1111111111111111101, 19'b1111111111111100101, 19'b0000000000000101101, 19'b1111111111110111000, 19'b0000000000001000100, 19'b1111111111101000101, 19'b0000000000000101001, 19'b1111111111111111111, 19'b0000000000001010000}, 
{19'b1111111111111101010, 19'b0000000000000000000, 19'b0000000000000101101, 19'b0000000000000000000, 19'b1111111111111100000, 19'b1111111111111111110, 19'b0000000000000110100, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000000000010, 19'b0000000000000000000, 19'b0000000000000001010, 19'b1111111111111001001, 19'b0000000000000000101, 19'b0000000000000111000, 19'b0000000000000010111, 19'b0000000000000110110, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000001000001, 19'b0000000000001111110, 19'b1111111111111001101, 19'b0000000000000000000, 19'b1111111111111111110, 19'b0000000000000000101, 19'b1111111111100010011, 19'b1111111111111111111, 19'b1111111111111011011, 19'b1111111111111111111, 19'b0000000000100100001, 19'b0000000000000000000, 19'b1111111111110010110}, 
{19'b1111111111111110010, 19'b1111111111111000010, 19'b1111111111111111011, 19'b0000000000000000011, 19'b0000000000000101110, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111111110100, 19'b0000000000000100100, 19'b1111111111111111011, 19'b0000000000000000000, 19'b0000000000000010000, 19'b0000000000010010111, 19'b1111111111111001011, 19'b0000000000000000110, 19'b1111111111001001101, 19'b1111111111111111010, 19'b1111111111111100001, 19'b0000000000000000100, 19'b1111111111111100110, 19'b0000000000000101111, 19'b1111111111110001101, 19'b0000000000000111010, 19'b0000000000000110101, 19'b1111111111111111001, 19'b1111111111010010011, 19'b1111111111110001010, 19'b1111111111111110100, 19'b1111111111111110110, 19'b0000000000011000111, 19'b1111111111111111101, 19'b0000000000001001110}, 
{19'b0000000000000011000, 19'b0000000000000000000, 19'b0000000000001011001, 19'b1111111111111000101, 19'b1111111111111011100, 19'b0000000000001111001, 19'b1111111111110101110, 19'b0000000000000011101, 19'b1111111111101100001, 19'b0000000000000000100, 19'b0000000000000001000, 19'b1111111111111010101, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111110011111, 19'b0000000000011011101, 19'b1111111111110000001, 19'b1111111111111111001, 19'b0000000000000111100, 19'b1111111111111111111, 19'b0000000000000100011, 19'b1111111111100001010, 19'b0000000000010100000, 19'b1111111111111111111, 19'b1111111111111000000, 19'b0000000000011111000, 19'b0000000000001001010, 19'b1111111111110101111, 19'b1111111111110111011, 19'b1111111111011101100, 19'b1111111111111111010, 19'b0000000000000001000}, 
{19'b1111111111111111111, 19'b0000000000000000011, 19'b1111111111111101110, 19'b1111111111101110110, 19'b1111111111111111111, 19'b1111111111100110111, 19'b0000000000000000000, 19'b0000000000010011011, 19'b0000000000001111101, 19'b0000000000000001001, 19'b0000000000000000000, 19'b1111111111111000111, 19'b0000000000010101010, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000011011110, 19'b0000000000000000000, 19'b1111111111111101011, 19'b1111111111111100101, 19'b1111111111101011011, 19'b0000000000001000011, 19'b0000000000000000000, 19'b0000000000000000000, 19'b0000000000000010000, 19'b1111111111111011011, 19'b1111111111100010100, 19'b0000000000010001101, 19'b1111111111100011100, 19'b0000000000000011010, 19'b1111111111111010111, 19'b0000000000000000000}, 
{19'b0000000000000011111, 19'b0000000000001011111, 19'b0000000000000000100, 19'b1111111111111111110, 19'b1111111111100010100, 19'b0000000000000000000, 19'b1111111111111111111, 19'b0000000000001111100, 19'b0000000000010001101, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000000000001, 19'b0000000000000000000, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111111111111, 19'b0000000000001010111, 19'b1111111111111001011, 19'b1111111111100100010, 19'b1111111111111101111, 19'b1111111111111001101, 19'b1111111111111001111, 19'b1111111111111011100, 19'b1111111111111111111, 19'b1111111111111011111, 19'b1111111111111110100, 19'b1111111111111111010, 19'b0000000000001001000, 19'b1111111111111111111, 19'b0000000000011101101}
};

localparam logic signed [18:0] bias [32] = '{
19'b0000000001011110010,  // 1.474280834197998
19'b0000000000101100010,  // 0.6914801001548767
19'b0000000001011100001,  // 1.4406442642211914
19'b0000000001011010000,  // 1.408045768737793
19'b0000000000111111001,  // 0.9864811301231384
19'b0000000000110111010,  // 0.8636202812194824
19'b1111111111011000100,  // -0.6153604388237
19'b0000000000011110111,  // 0.4839226007461548
19'b0000000000011111000,  // 0.4862793982028961
19'b0000000000010111110,  // 0.37162142992019653
19'b0000000000011101011,  // 0.45989668369293213
19'b0000000001010011001,  // 1.2998151779174805
19'b1111111110111110111,  // -1.016528844833374
19'b1111111111101001011,  // -0.35249894857406616
19'b0000000000011100100,  // 0.44582197070121765
19'b1111111111111000110,  // -0.1119980737566948
19'b1111111111111011101,  // -0.06717441976070404
19'b0000000000000000010,  // 0.00487547367811203
19'b0000000000001100011,  // 0.1946917623281479
19'b1111111111001110000,  // -0.7796769738197327
19'b0000000000101110101,  // 0.7287401556968689
19'b0000000001101101110,  // 1.714877724647522
19'b1111111110011001110,  // -1.5971007347106934
19'b0000000000000100101,  // 0.07393483817577362
19'b0000000000010100101,  // 0.3225609362125397
19'b0000000000110110000,  // 0.8453295230865479
19'b0000000000111001100,  // 0.898597240447998
19'b0000000000010000010,  // 0.2548799514770508
19'b0000000000111110010,  // 0.9735668301582336
19'b0000000001001000000,  // 1.1261906623840332
19'b0000000000011100101,  // 0.44768181443214417
19'b1111111101101000011   // -2.3676068782806396
};
endpackage