// Width: 12
// NFRAC: 6
package dense_4_12_6;

localparam logic signed [11:0] weights [32][5] = '{ 
{12'b111111111111, 12'b000000010100, 12'b111111101100, 12'b000000000100, 12'b111111111001}, 
{12'b111111011100, 12'b111111111100, 12'b000000011101, 12'b111111111111, 12'b000000000001}, 
{12'b000000010111, 12'b000000001101, 12'b111111111110, 12'b111111100110, 12'b111111110010}, 
{12'b111111100111, 12'b111111101000, 12'b111111111000, 12'b000000010011, 12'b000000001111}, 
{12'b000000000111, 12'b000000001000, 12'b000000001010, 12'b111111111110, 12'b111110111111}, 
{12'b000000010100, 12'b111111100110, 12'b000000001011, 12'b111111110101, 12'b111111110101}, 
{12'b111111100110, 12'b000000000010, 12'b111111111111, 12'b000000001011, 12'b000000000100}, 
{12'b111111111111, 12'b000000010010, 12'b111111100110, 12'b000000001010, 12'b000000001000}, 
{12'b000000001010, 12'b111111110101, 12'b000000000000, 12'b111111100010, 12'b111111110000}, 
{12'b111111111111, 12'b111111101110, 12'b000000001011, 12'b000000011011, 12'b000000000000}, 
{12'b111111110111, 12'b111111110110, 12'b000000000000, 12'b000000100101, 12'b111111101110}, 
{12'b000000001010, 12'b000000001110, 12'b111111101010, 12'b111111111110, 12'b000000000111}, 
{12'b000000000000, 12'b000000001010, 12'b000000000000, 12'b111111110010, 12'b111111011000}, 
{12'b000000001011, 12'b000000000100, 12'b000000011010, 12'b111111111011, 12'b111111100100}, 
{12'b000000000101, 12'b111111111100, 12'b111111101000, 12'b111111111101, 12'b000000100010}, 
{12'b111111100001, 12'b111111110000, 12'b111111110001, 12'b000000011001, 12'b000000000010}, 
{12'b000000010110, 12'b111111110101, 12'b111111110111, 12'b111111110001, 12'b111111111100}, 
{12'b000000001100, 12'b111111111101, 12'b111111100101, 12'b111111111110, 12'b000000000100}, 
{12'b000000010000, 12'b000000000010, 12'b111111110010, 12'b000000000000, 12'b111111100111}, 
{12'b000000001110, 12'b111111111010, 12'b111111110010, 12'b000000001101, 12'b000000000110}, 
{12'b000000000100, 12'b111111111110, 12'b000000010011, 12'b111111100100, 12'b111111111110}, 
{12'b000000000000, 12'b000000000111, 12'b000000011111, 12'b111111011110, 12'b111111011000}, 
{12'b111111111001, 12'b000000000111, 12'b000000001011, 12'b111111101001, 12'b000000100001}, 
{12'b111111111111, 12'b000000001010, 12'b000000010010, 12'b000000000010, 12'b111111011011}, 
{12'b111111110101, 12'b000000010111, 12'b111111110001, 12'b000000000000, 12'b000000011000}, 
{12'b000000000001, 12'b000000010001, 12'b000000000001, 12'b111111010000, 12'b000000100011}, 
{12'b111111100010, 12'b111111110000, 12'b000000001101, 12'b000000001111, 12'b000000001100}, 
{12'b000000000000, 12'b000000001111, 12'b111111111101, 12'b111111110110, 12'b000000000010}, 
{12'b111111111001, 12'b000000001111, 12'b111111011111, 12'b000000001000, 12'b111111110101}, 
{12'b111111111110, 12'b000000001001, 12'b111111110101, 12'b111111100110, 12'b000000100101}, 
{12'b000000011100, 12'b000000000100, 12'b000000010100, 12'b111111011010, 12'b111111101011}, 
{12'b111111111100, 12'b111111100111, 12'b000000010111, 12'b000000000100, 12'b000000001000}
};

localparam logic signed [11:0] bias [5] = '{
12'b111111111100,  // -0.06223141402006149
12'b111111111011,  // -0.06270556896924973
12'b111111111011,  // -0.07014333456754684
12'b000000000101,  // 0.0820775106549263
12'b000000001101   // 0.2155742198228836
};
endpackage