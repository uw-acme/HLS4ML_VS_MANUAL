// Width: 9
// NFRAC: 4
package dense_2_9_5;

localparam logic signed [8:0] weights [64][32] = '{ 
{9'b000000100, 9'b000000000, 9'b111111100, 9'b111111111, 9'b000000100, 9'b000000000, 9'b111111101, 9'b111111111, 9'b111111011, 9'b000000001, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111100, 9'b111111111, 9'b111111011, 9'b000000000, 9'b111111111, 9'b111111100, 9'b111111101, 9'b000000000, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000001, 9'b000000110, 9'b000000010, 9'b111111111, 9'b000000000, 9'b111111001, 9'b000000000}, 
{9'b111111110, 9'b111111101, 9'b111111101, 9'b111111111, 9'b111111111, 9'b000000000, 9'b111111100, 9'b000000000, 9'b000000000, 9'b111111110, 9'b000000010, 9'b111111111, 9'b111111111, 9'b111111100, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111100, 9'b000000010, 9'b000000011, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000000, 9'b111111110, 9'b000000100, 9'b000000011, 9'b000000000, 9'b000000000, 9'b111111000, 9'b000000000, 9'b000000000}, 
{9'b000000001, 9'b111111110, 9'b111111101, 9'b111111111, 9'b111111110, 9'b111111110, 9'b111111101, 9'b000000000, 9'b111111101, 9'b000000000, 9'b000000000, 9'b111111110, 9'b000000001, 9'b111111110, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000001, 9'b000000000, 9'b000000011, 9'b000000000, 9'b111111110, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000011, 9'b000000010, 9'b000000001, 9'b111111111, 9'b111111101, 9'b111111111, 9'b000000001}, 
{9'b000000010, 9'b000000000, 9'b000000000, 9'b111111111, 9'b111110111, 9'b000000000, 9'b000000000, 9'b000000011, 9'b000000011, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000011, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111101, 9'b111111111, 9'b000000000, 9'b111111110, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000001, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111100, 9'b000000100}, 
{9'b111110101, 9'b111111111, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111111, 9'b111111101, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000011, 9'b000000000, 9'b000000101, 9'b111111111, 9'b000000011, 9'b111111001, 9'b000000000, 9'b111111110, 9'b000000010, 9'b000000100, 9'b000000000, 9'b000000000, 9'b000000010, 9'b000000011, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000011}, 
{9'b000000000, 9'b111111111, 9'b000000010, 9'b111110101, 9'b111101001, 9'b111111010, 9'b000000101, 9'b111110110, 9'b111111111, 9'b111110101, 9'b111110111, 9'b111111010, 9'b000000101, 9'b111111111, 9'b111111111, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111101, 9'b111111111, 9'b111111000, 9'b000000000, 9'b000000010, 9'b111111111, 9'b000000000, 9'b000000100, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000011, 9'b111111111, 9'b000000011}, 
{9'b111111111, 9'b111111101, 9'b111111100, 9'b111111111, 9'b111111011, 9'b000000001, 9'b111111101, 9'b111111101, 9'b111111001, 9'b000000000, 9'b111111111, 9'b111111101, 9'b000000001, 9'b111111111, 9'b111111111, 9'b111110111, 9'b111111111, 9'b000000001, 9'b000000011, 9'b111111101, 9'b111111101, 9'b111111110, 9'b111111111, 9'b000000000, 9'b111111111, 9'b111110101, 9'b111111011, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111111}, 
{9'b111111101, 9'b111111110, 9'b111111110, 9'b111111100, 9'b111111110, 9'b111111111, 9'b000000001, 9'b111111110, 9'b000000011, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000011, 9'b000000000, 9'b111111111, 9'b111111110, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111101, 9'b000000000, 9'b111111111, 9'b111111110, 9'b111111111, 9'b000000000, 9'b111111111}, 
{9'b111111000, 9'b111111111, 9'b111111001, 9'b000000001, 9'b000000111, 9'b111111111, 9'b111111111, 9'b000000011, 9'b111111000, 9'b111111111, 9'b000000000, 9'b111111100, 9'b111111111, 9'b000000001, 9'b111111100, 9'b000001100, 9'b111111111, 9'b000000000, 9'b000000011, 9'b000000011, 9'b000000000, 9'b111111010, 9'b000000000, 9'b000000110, 9'b111111101, 9'b000001011, 9'b111111101, 9'b111111100, 9'b111111000, 9'b111111000, 9'b000000000, 9'b000000000}, 
{9'b000000000, 9'b111111111, 9'b111111110, 9'b000000000, 9'b000000100, 9'b111111111, 9'b111111110, 9'b000000001, 9'b000000001, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111110, 9'b111111111, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000000, 9'b000000001, 9'b000000000, 9'b111111111, 9'b000000000, 9'b000000000, 9'b000000000, 9'b111111101, 9'b000000001, 9'b000000011, 9'b111111111, 9'b000000000, 9'b000000000, 9'b000000001}, 
{9'b000000001, 9'b000000000, 9'b111111110, 9'b111111011, 9'b111110011, 9'b000000010, 9'b000000000, 9'b111110010, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000000, 9'b000000000, 9'b111111111, 9'b111111001, 9'b111111111, 9'b000000011, 9'b000000010, 9'b000000011, 9'b111111000, 9'b111111010, 9'b000000001, 9'b111111111, 9'b111111111, 9'b000000101, 9'b111111110, 9'b111111111, 9'b111111111, 9'b000000011, 9'b111111111, 9'b000000000}, 
{9'b111111100, 9'b111111000, 9'b000000000, 9'b111111111, 9'b000000101, 9'b111111011, 9'b111111100, 9'b000000001, 9'b111111111, 9'b000000010, 9'b000000001, 9'b111111110, 9'b000000000, 9'b000000000, 9'b111111111, 9'b111111011, 9'b000000010, 9'b000000000, 9'b000000100, 9'b000000001, 9'b000000000, 9'b111111111, 9'b000000010, 9'b111111110, 9'b111111011, 9'b111111111, 9'b000000010, 9'b111111111, 9'b000000000, 9'b111111110, 9'b000000010, 9'b000000100}, 
{9'b000000000, 9'b000000000, 9'b000000011, 9'b000000000, 9'b111111111, 9'b000000010, 9'b000000001, 9'b111111111, 9'b000000000, 9'b111111101, 9'b111111111, 9'b111111101, 9'b111111111, 9'b000000000, 9'b111111110, 9'b000001101, 9'b000000000, 9'b111111110, 9'b111111100, 9'b111111111, 9'b000000011, 9'b000000010, 9'b000000000, 9'b111111111, 9'b000000011, 9'b000000100, 9'b000000111, 9'b000000000, 9'b000000000, 9'b000000000, 9'b111111111, 9'b111111110}, 
{9'b111111101, 9'b000000000, 9'b000000000, 9'b111111100, 9'b111111011, 9'b000000111, 9'b000000000, 9'b000000000, 9'b111111101, 9'b111111110, 9'b000000010, 9'b000000001, 9'b000000000, 9'b111111110, 9'b000000100, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000001, 9'b000000000, 9'b000000001, 9'b111111111, 9'b000000000, 9'b000001010, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111110, 9'b111111111, 9'b000000010}, 
{9'b000000000, 9'b000000001, 9'b000000101, 9'b111111111, 9'b000000001, 9'b000000101, 9'b000000000, 9'b111111111, 9'b000000001, 9'b111111110, 9'b111111111, 9'b111111110, 9'b000000000, 9'b000000110, 9'b111111111, 9'b000000000, 9'b000000011, 9'b000000000, 9'b000000000, 9'b111111010, 9'b111111100, 9'b111111111, 9'b111111111, 9'b111111101, 9'b111111111, 9'b111111110, 9'b111111100, 9'b111111100, 9'b000000000, 9'b000000001, 9'b111111001, 9'b000000000}, 
{9'b111111011, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000010, 9'b111111110, 9'b000000100, 9'b111111010, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000000, 9'b000000000, 9'b111111111, 9'b111111110, 9'b000000001, 9'b000000010, 9'b111111111, 9'b111111011, 9'b111111111, 9'b000000001, 9'b000000001, 9'b000000000, 9'b000000000, 9'b000000001, 9'b111111100, 9'b000000000, 9'b111111111, 9'b000000000, 9'b000000000, 9'b111111101}, 
{9'b111111010, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000001, 9'b000000000, 9'b000000000, 9'b000000000, 9'b000000001, 9'b000000001, 9'b000000010, 9'b000000000, 9'b111111110, 9'b000000000, 9'b000000110, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000001, 9'b000000010, 9'b000000000, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000000, 9'b111111110, 9'b111111101, 9'b000000011, 9'b111111111, 9'b000000000, 9'b111111100}, 
{9'b000000000, 9'b111111111, 9'b000000000, 9'b000000000, 9'b000001110, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000001, 9'b111111110, 9'b000000000, 9'b000000000, 9'b000000000, 9'b000000010, 9'b000000000, 9'b111111101, 9'b111111111, 9'b111111110, 9'b000000101, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000000, 9'b000000001, 9'b000000000, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000000}, 
{9'b111111111, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111111, 9'b111111110, 9'b111111111, 9'b000000100, 9'b000000000, 9'b000000001, 9'b111111111, 9'b000000001, 9'b111111111, 9'b111111101, 9'b111111100, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000001, 9'b000000000, 9'b111111101, 9'b000000001, 9'b111111101, 9'b000000000, 9'b000000000, 9'b111111101, 9'b000000000, 9'b000000000, 9'b111111111}, 
{9'b111111111, 9'b111111110, 9'b000000000, 9'b111111111, 9'b000000011, 9'b111111111, 9'b111111111, 9'b000000001, 9'b111111001, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000101, 9'b000000011, 9'b111111110, 9'b111111111, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000000, 9'b000000000, 9'b111111101, 9'b111111110, 9'b000000010, 9'b000000000, 9'b111111101, 9'b000000000, 9'b111111110, 9'b111111111, 9'b000000010, 9'b000000000, 9'b111111100}, 
{9'b000001010, 9'b000000101, 9'b111111100, 9'b000000000, 9'b111111010, 9'b000000000, 9'b000000011, 9'b000000000, 9'b000000011, 9'b111111111, 9'b111111101, 9'b111111110, 9'b000000010, 9'b000000000, 9'b111111110, 9'b000000010, 9'b000001000, 9'b111111101, 9'b111111011, 9'b000000000, 9'b111111111, 9'b111111101, 9'b111111111, 9'b111111111, 9'b000000001, 9'b111111010, 9'b000000001, 9'b111111111, 9'b000000000, 9'b000000001, 9'b111111111, 9'b000000000}, 
{9'b111111110, 9'b111111100, 9'b111111111, 9'b111111101, 9'b111111111, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111100, 9'b000000001, 9'b000000001, 9'b111111110, 9'b000000111, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000000, 9'b000000101, 9'b111111000, 9'b111111110, 9'b111111111, 9'b111111111, 9'b000000011, 9'b111111111, 9'b000000000, 9'b000000111, 9'b111110111, 9'b111111010, 9'b000000000}, 
{9'b000000000, 9'b111111111, 9'b111111111, 9'b000000000, 9'b111110100, 9'b111110110, 9'b000000000, 9'b111111111, 9'b111111011, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111110, 9'b111111101, 9'b000000100, 9'b000000000, 9'b000000000, 9'b111111111, 9'b111111110, 9'b000000000, 9'b111111110, 9'b000000011, 9'b111110110, 9'b000000011, 9'b111111111, 9'b111111111, 9'b000000011, 9'b111111111, 9'b000000011}, 
{9'b111111111, 9'b000000000, 9'b111111111, 9'b000000001, 9'b000000000, 9'b111111010, 9'b000000000, 9'b000000001, 9'b000001001, 9'b111111111, 9'b000000000, 9'b000000000, 9'b000000101, 9'b111111111, 9'b000000000, 9'b000000001, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111011, 9'b000000000, 9'b000000001, 9'b000000000, 9'b111111111, 9'b000000011, 9'b000000000, 9'b000000010, 9'b111111001, 9'b000000001, 9'b000000110, 9'b000000000}, 
{9'b111111010, 9'b000000011, 9'b111111011, 9'b000000001, 9'b111111110, 9'b000000000, 9'b000000111, 9'b111111100, 9'b111111011, 9'b000000010, 9'b111111100, 9'b111111111, 9'b111111111, 9'b000000101, 9'b111111111, 9'b111111011, 9'b111111111, 9'b000000111, 9'b111111000, 9'b111111111, 9'b000000101, 9'b111111010, 9'b000000000, 9'b111111111, 9'b000000100, 9'b111110111, 9'b111111010, 9'b111111100, 9'b111111111, 9'b000000001, 9'b000000000, 9'b000000010}, 
{9'b111111110, 9'b000000000, 9'b111111111, 9'b000000010, 9'b111111111, 9'b000000011, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000001000, 9'b000000000, 9'b000000011, 9'b000000000, 9'b111111100, 9'b111111110, 9'b111111111, 9'b111111111, 9'b000000000, 9'b111111111, 9'b111111101, 9'b111111111, 9'b000000100, 9'b000000100, 9'b111111111, 9'b111111111, 9'b000000000, 9'b111111111, 9'b111111110}, 
{9'b111111110, 9'b000000000, 9'b000000100, 9'b000000000, 9'b000000000, 9'b111111110, 9'b000000000, 9'b111110010, 9'b000000011, 9'b000000000, 9'b000000000, 9'b111111010, 9'b000000000, 9'b111111101, 9'b111111111, 9'b000000000, 9'b000000000, 9'b000000000, 9'b000000001, 9'b000000000, 9'b111111111, 9'b000000101, 9'b000000110, 9'b111111100, 9'b111111101, 9'b000000011, 9'b111111011, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000010}, 
{9'b111111110, 9'b111111111, 9'b111111100, 9'b111111100, 9'b111111111, 9'b111111101, 9'b000000000, 9'b000000001, 9'b111111100, 9'b111111110, 9'b111111111, 9'b000000000, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000001, 9'b000000011, 9'b000000010, 9'b111111101, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000000, 9'b111111110, 9'b000000001, 9'b111111110, 9'b000000000, 9'b111111111, 9'b111111011, 9'b111111111, 9'b000000011}, 
{9'b111111111, 9'b111111110, 9'b000000001, 9'b000000100, 9'b000000001, 9'b000000001, 9'b000000000, 9'b111111100, 9'b111111100, 9'b000000001, 9'b000000000, 9'b000000000, 9'b000000000, 9'b000000000, 9'b000000011, 9'b000000000, 9'b111111111, 9'b000000001, 9'b111111111, 9'b111111111, 9'b000000001, 9'b111111110, 9'b111111111, 9'b000000010, 9'b000000000, 9'b111111110, 9'b111111100, 9'b111111111, 9'b111111011, 9'b000000000, 9'b000000001, 9'b000000000}, 
{9'b111111111, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111101, 9'b111111101, 9'b000000001, 9'b000000000, 9'b111111101, 9'b000000010, 9'b111111111, 9'b111111111, 9'b111111110, 9'b000000000, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111110, 9'b000000000, 9'b111111101, 9'b000000001, 9'b111111100, 9'b000000000, 9'b000000000, 9'b000000001, 9'b000000000, 9'b000000000, 9'b000000100, 9'b000000000, 9'b000000000, 9'b000000001}, 
{9'b111111111, 9'b000000100, 9'b111111111, 9'b111111111, 9'b111111100, 9'b111111110, 9'b000000110, 9'b111110100, 9'b111111010, 9'b111111100, 9'b111111100, 9'b111111011, 9'b111111111, 9'b000000111, 9'b111111111, 9'b000000000, 9'b111111100, 9'b000000111, 9'b111111001, 9'b000000000, 9'b111111111, 9'b111111010, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111111, 9'b111111101, 9'b111111111, 9'b000000010, 9'b000000000, 9'b111111110, 9'b000000000}, 
{9'b000000101, 9'b111111110, 9'b000000010, 9'b111111111, 9'b000000001, 9'b111111111, 9'b111111111, 9'b111111110, 9'b000000000, 9'b000000001, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000011, 9'b000000000, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000000, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111011, 9'b111111111, 9'b000000000, 9'b111111110, 9'b111111101, 9'b111111111, 9'b111111111, 9'b000001000, 9'b111111011, 9'b111111110}, 
{9'b111111111, 9'b111111110, 9'b111111110, 9'b000000000, 9'b000000010, 9'b111111101, 9'b111111111, 9'b111111100, 9'b000000000, 9'b000000010, 9'b111111100, 9'b111111011, 9'b000000000, 9'b111110101, 9'b111111110, 9'b111111110, 9'b111111100, 9'b111111111, 9'b000000010, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000000, 9'b111111111, 9'b111110011, 9'b111110111, 9'b111111011, 9'b000000000, 9'b000000011, 9'b111111111, 9'b000000011}, 
{9'b111111110, 9'b111111100, 9'b000000010, 9'b000000001, 9'b000000000, 9'b111111110, 9'b111111111, 9'b000000001, 9'b000001000, 9'b111111101, 9'b111111111, 9'b111111111, 9'b000000001, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111110, 9'b111111111, 9'b000000000, 9'b000000011, 9'b111111101, 9'b111111111, 9'b000000010, 9'b111111111, 9'b000000000, 9'b000001000, 9'b000000101, 9'b000000000, 9'b000000000, 9'b111111001, 9'b111111110, 9'b111111111}, 
{9'b000000000, 9'b000000000, 9'b111111111, 9'b000000000, 9'b000000011, 9'b111111000, 9'b000000000, 9'b111111110, 9'b000000010, 9'b000000000, 9'b111111111, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111110, 9'b000000100, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111010, 9'b000000000, 9'b000000010, 9'b111111111, 9'b000000001, 9'b111111111, 9'b000000001}, 
{9'b111111100, 9'b000000000, 9'b111111000, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111110, 9'b111111111, 9'b111111110, 9'b000000000, 9'b000000000, 9'b111111101, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000001, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000100, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000101, 9'b000000011, 9'b000000000, 9'b111111110, 9'b111111111, 9'b000000001, 9'b000000000}, 
{9'b000000000, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111000, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111101, 9'b111111111, 9'b000000000, 9'b111111101, 9'b000000000, 9'b000000000, 9'b000000000, 9'b000000000, 9'b111111010, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000010, 9'b111111111, 9'b000000000, 9'b000000111, 9'b000000101, 9'b000000000, 9'b000000000, 9'b111111100, 9'b000000000, 9'b111111111}, 
{9'b000000001, 9'b000000000, 9'b000000100, 9'b111111100, 9'b000000010, 9'b000000001, 9'b000000000, 9'b000000011, 9'b000000000, 9'b111111111, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000001, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000001, 9'b000000000, 9'b111110110, 9'b111111110, 9'b000000001, 9'b111111111, 9'b111110111, 9'b111111101, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000000, 9'b111111111}, 
{9'b000000000, 9'b111111111, 9'b111111110, 9'b111111101, 9'b000000000, 9'b000000000, 9'b000000001, 9'b111111111, 9'b000000011, 9'b111111111, 9'b000000000, 9'b111111010, 9'b111111111, 9'b000000010, 9'b111111111, 9'b111111011, 9'b000000000, 9'b111111111, 9'b000000100, 9'b111111111, 9'b111111001, 9'b111111111, 9'b000000100, 9'b111111111, 9'b111111111, 9'b000000010, 9'b111111110, 9'b000000001, 9'b000000000, 9'b111111100, 9'b000000000, 9'b000000000}, 
{9'b111111100, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000111, 9'b111111110, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000001, 9'b000000010, 9'b111111111, 9'b000000011, 9'b000000000, 9'b111111111, 9'b111111011, 9'b111111111, 9'b000000000, 9'b111111110, 9'b000000000, 9'b000000000, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111100, 9'b111111011, 9'b000000000, 9'b111111110, 9'b000000000, 9'b111111111, 9'b000000001}, 
{9'b111111001, 9'b111111101, 9'b111111101, 9'b000000000, 9'b000001001, 9'b111111100, 9'b000000000, 9'b111111111, 9'b111111001, 9'b000000010, 9'b111111111, 9'b000001001, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000111, 9'b000000000, 9'b111111111, 9'b000000001, 9'b111111111, 9'b111111111, 9'b111111110, 9'b111111111, 9'b111111000, 9'b111111101, 9'b111111111, 9'b111111111, 9'b111111111}, 
{9'b000000011, 9'b111110011, 9'b111110100, 9'b111111101, 9'b000001010, 9'b111111111, 9'b111111010, 9'b000000100, 9'b000000000, 9'b000000000, 9'b000000011, 9'b111111011, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111110, 9'b111110001, 9'b000000010, 9'b000000101, 9'b000000100, 9'b000000000, 9'b000000000, 9'b111111001, 9'b111110101, 9'b111111111, 9'b111111011, 9'b111111000, 9'b111111100, 9'b111110001, 9'b000000110, 9'b000000110}, 
{9'b000000000, 9'b000000000, 9'b000000000, 9'b000000000, 9'b000000100, 9'b111111101, 9'b000000000, 9'b000000001, 9'b111111010, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000011, 9'b000000000, 9'b000000000, 9'b000000000, 9'b000000101, 9'b111111100, 9'b000000000, 9'b111111101, 9'b111111111, 9'b000000101, 9'b000000000, 9'b111111111, 9'b111110111, 9'b111111111, 9'b111111101, 9'b111111111, 9'b000000000, 9'b000000010, 9'b000000001}, 
{9'b111111111, 9'b000000010, 9'b111111011, 9'b000000000, 9'b000000011, 9'b111111111, 9'b111111111, 9'b000000010, 9'b000000000, 9'b111111111, 9'b111111110, 9'b000000000, 9'b000000000, 9'b111111111, 9'b111111110, 9'b111111110, 9'b111111111, 9'b111111110, 9'b111111110, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111110, 9'b000000110, 9'b000000000, 9'b111111010, 9'b111111111, 9'b000000001, 9'b000000000, 9'b000000000, 9'b000000100, 9'b111111111}, 
{9'b111111111, 9'b000000000, 9'b111111111, 9'b111111101, 9'b111110010, 9'b000000000, 9'b000000000, 9'b111111111, 9'b111110110, 9'b000000001, 9'b111111110, 9'b111111111, 9'b000000000, 9'b111111010, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000000, 9'b000000000, 9'b000000101, 9'b111111110, 9'b111111011, 9'b000000000, 9'b111111011, 9'b111111110, 9'b111111100, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111000, 9'b111111111, 9'b000000011}, 
{9'b000000001, 9'b000000011, 9'b111111111, 9'b000000010, 9'b111111100, 9'b111111110, 9'b000000001, 9'b000000001, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111010, 9'b111111111, 9'b000000010, 9'b111111110, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000011, 9'b111111010, 9'b000000100, 9'b000000000, 9'b000000000, 9'b000000011, 9'b000000000, 9'b111111111, 9'b111111001, 9'b111111110, 9'b111111101, 9'b000000010}, 
{9'b000000000, 9'b000000000, 9'b111111010, 9'b111111111, 9'b000000011, 9'b111111101, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000000, 9'b000000000, 9'b111111100, 9'b000000001, 9'b000000000, 9'b000000000, 9'b000000000, 9'b111111111, 9'b111111101, 9'b000000000, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000100, 9'b111111111, 9'b000000000, 9'b111111011, 9'b111111010, 9'b000000011, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000100}, 
{9'b111111010, 9'b111111111, 9'b111111100, 9'b000000000, 9'b111111010, 9'b000000000, 9'b111111111, 9'b111111110, 9'b111110111, 9'b111111111, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111101, 9'b111111110, 9'b000000001, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000101, 9'b111111111, 9'b000000010, 9'b000000001, 9'b111111101, 9'b000000011, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000001001}, 
{9'b111111010, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000011, 9'b111111011, 9'b111111111, 9'b000000100, 9'b000000010, 9'b000000000, 9'b111111111, 9'b111111110, 9'b111111110, 9'b111111110, 9'b111111111, 9'b000000001, 9'b111111111, 9'b000000000, 9'b000000010, 9'b000000000, 9'b000000000, 9'b000000000, 9'b000000100, 9'b000000000, 9'b000000000, 9'b111111110, 9'b111111111, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000001}, 
{9'b111111111, 9'b000000000, 9'b111111100, 9'b111111110, 9'b000000100, 9'b111111111, 9'b111111110, 9'b000000011, 9'b111111111, 9'b000000100, 9'b000000001, 9'b111111110, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111110, 9'b111111011, 9'b000000100, 9'b000000010, 9'b000001010, 9'b000000011, 9'b000000011, 9'b111111111, 9'b000000000, 9'b000000000, 9'b000000000, 9'b000000001, 9'b111111001, 9'b111111111, 9'b111111111, 9'b111111111}, 
{9'b000000000, 9'b111111110, 9'b111111110, 9'b000000000, 9'b111111100, 9'b000000000, 9'b000000011, 9'b000000001, 9'b000000000, 9'b111111110, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000011, 9'b111111111, 9'b111111111, 9'b111111011, 9'b000000000, 9'b111111100, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000000, 9'b000000000, 9'b000000000, 9'b000000010, 9'b111111110, 9'b111111111, 9'b111111000, 9'b000000001}, 
{9'b000000111, 9'b111111111, 9'b000000001, 9'b111111110, 9'b111111110, 9'b000000000, 9'b000000010, 9'b000000000, 9'b000001000, 9'b000000000, 9'b111111111, 9'b000000000, 9'b000000001, 9'b111111111, 9'b000000000, 9'b000000001, 9'b111111111, 9'b111111000, 9'b111111111, 9'b111111111, 9'b000000001, 9'b000000000, 9'b111111111, 9'b000000001, 9'b000000000, 9'b111111011, 9'b111111110, 9'b000000010, 9'b111111111, 9'b000000100, 9'b111111111, 9'b111111101}, 
{9'b000000000, 9'b000000001, 9'b111111111, 9'b111111111, 9'b111111010, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000010, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000101, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000010, 9'b000000000, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000000, 9'b000000000, 9'b000000000, 9'b000000001}, 
{9'b111111011, 9'b000000010, 9'b000000000, 9'b111111110, 9'b111111001, 9'b111111111, 9'b000000001, 9'b111111001, 9'b000001000, 9'b000000001, 9'b000000000, 9'b000000001, 9'b000000000, 9'b000000000, 9'b000000110, 9'b111111110, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111001, 9'b000000000, 9'b000000010, 9'b000000000, 9'b000000000, 9'b111110101, 9'b111111010, 9'b111111100, 9'b000000000, 9'b111111111, 9'b000000101, 9'b111111100}, 
{9'b111111111, 9'b111111100, 9'b111111110, 9'b111111001, 9'b111111011, 9'b000000101, 9'b000000100, 9'b111111101, 9'b000000000, 9'b111111111, 9'b111111110, 9'b111111011, 9'b000000001, 9'b111111011, 9'b000000011, 9'b111111111, 9'b000000101, 9'b111111111, 9'b111111111, 9'b111111101, 9'b111111111, 9'b111111110, 9'b111111011, 9'b000000001, 9'b111111111, 9'b111111111, 9'b111111100, 9'b000000101, 9'b000000100, 9'b111111110, 9'b111110101, 9'b000000010}, 
{9'b000000000, 9'b111111111, 9'b111111111, 9'b111111110, 9'b000000000, 9'b000000000, 9'b000000001, 9'b000000000, 9'b000000001, 9'b111111111, 9'b000000000, 9'b000000001, 9'b000000000, 9'b000000000, 9'b111111101, 9'b111111110, 9'b000000000, 9'b000000010, 9'b000000000, 9'b000000010, 9'b111111111, 9'b111111101, 9'b111111111, 9'b000000001, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000001, 9'b000000000, 9'b000000001, 9'b111111001, 9'b111111111}, 
{9'b000000100, 9'b111111111, 9'b000000010, 9'b111111011, 9'b111111100, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000000, 9'b111111101, 9'b000000000, 9'b000000000, 9'b000000000, 9'b000000000, 9'b111111101, 9'b000000010, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000001, 9'b111111100, 9'b000000001, 9'b000000010, 9'b000000010, 9'b111111111, 9'b000001000, 9'b111111101, 9'b000000101, 9'b111111111, 9'b111111010, 9'b111111101, 9'b000000010}, 
{9'b111110111, 9'b111111111, 9'b111111101, 9'b111111111, 9'b000000100, 9'b111111101, 9'b111111111, 9'b000000011, 9'b000000001, 9'b111111100, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000010, 9'b111111100, 9'b111111111, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000000, 9'b111111100, 9'b111111111, 9'b000000000, 9'b111111010, 9'b000000001, 9'b000001001, 9'b000000101, 9'b111111111, 9'b111111101, 9'b111111000, 9'b000000000, 9'b111111111}, 
{9'b000000000, 9'b000000011, 9'b000000000, 9'b111111101, 9'b000000000, 9'b111111111, 9'b000000000, 9'b000000011, 9'b000000011, 9'b111111101, 9'b000000010, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111101, 9'b000000100, 9'b111111111, 9'b111111010, 9'b000000001, 9'b111111111, 9'b111111111, 9'b000000001, 9'b111111110, 9'b111111111, 9'b111111111, 9'b000000001, 9'b111111101, 9'b000000010, 9'b111111010, 9'b000000001, 9'b111111111, 9'b000000010}, 
{9'b111111111, 9'b000000000, 9'b000000001, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000001, 9'b111111111, 9'b000000000, 9'b000000000, 9'b000000000, 9'b000000000, 9'b111111110, 9'b000000000, 9'b000000001, 9'b000000000, 9'b000000001, 9'b111111111, 9'b111111111, 9'b000000010, 9'b000000011, 9'b111111110, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111000, 9'b111111111, 9'b111111110, 9'b111111111, 9'b000001001, 9'b000000000, 9'b111111100}, 
{9'b111111111, 9'b111111110, 9'b111111111, 9'b000000000, 9'b000000001, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000001, 9'b111111111, 9'b000000000, 9'b000000000, 9'b000000100, 9'b111111110, 9'b000000000, 9'b111110010, 9'b111111111, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000001, 9'b111111100, 9'b000000001, 9'b000000001, 9'b111111111, 9'b111110100, 9'b111111100, 9'b111111111, 9'b111111111, 9'b000000110, 9'b111111111, 9'b000000010}, 
{9'b000000000, 9'b000000000, 9'b000000010, 9'b111111110, 9'b111111110, 9'b000000011, 9'b111111101, 9'b000000000, 9'b111111011, 9'b000000000, 9'b000000000, 9'b111111110, 9'b000000000, 9'b000000000, 9'b111111100, 9'b000000110, 9'b111111100, 9'b111111111, 9'b000000001, 9'b111111111, 9'b000000001, 9'b111111000, 9'b000000101, 9'b111111111, 9'b111111110, 9'b000000111, 9'b000000010, 9'b111111101, 9'b111111101, 9'b111110111, 9'b111111111, 9'b000000000}, 
{9'b111111111, 9'b000000000, 9'b111111111, 9'b111111011, 9'b111111111, 9'b111111001, 9'b000000000, 9'b000000100, 9'b000000011, 9'b000000000, 9'b000000000, 9'b111111110, 9'b000000101, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000110, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111010, 9'b000000010, 9'b000000000, 9'b000000000, 9'b000000000, 9'b111111110, 9'b111111000, 9'b000000100, 9'b111111000, 9'b000000000, 9'b111111110, 9'b000000000}, 
{9'b000000000, 9'b000000010, 9'b000000000, 9'b111111111, 9'b111111000, 9'b000000000, 9'b111111111, 9'b000000011, 9'b000000100, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000000, 9'b000000000, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000010, 9'b111111110, 9'b111111001, 9'b111111111, 9'b111111110, 9'b111111110, 9'b111111110, 9'b111111111, 9'b111111110, 9'b111111111, 9'b111111111, 9'b000000010, 9'b111111111, 9'b000000111}
};

localparam logic signed [8:0] bias [32] = '{
9'b000010111,  // 1.474280834197998
9'b000001011,  // 0.6914801001548767
9'b000010111,  // 1.4406442642211914
9'b000010110,  // 1.408045768737793
9'b000001111,  // 0.9864811301231384
9'b000001101,  // 0.8636202812194824
9'b111110110,  // -0.6153604388237
9'b000000111,  // 0.4839226007461548
9'b000000111,  // 0.4862793982028961
9'b000000101,  // 0.37162142992019653
9'b000000111,  // 0.45989668369293213
9'b000010100,  // 1.2998151779174805
9'b111101111,  // -1.016528844833374
9'b111111010,  // -0.35249894857406616
9'b000000111,  // 0.44582197070121765
9'b111111110,  // -0.1119980737566948
9'b111111110,  // -0.06717441976070404
9'b000000000,  // 0.00487547367811203
9'b000000011,  // 0.1946917623281479
9'b111110011,  // -0.7796769738197327
9'b000001011,  // 0.7287401556968689
9'b000011011,  // 1.714877724647522
9'b111100110,  // -1.5971007347106934
9'b000000001,  // 0.07393483817577362
9'b000000101,  // 0.3225609362125397
9'b000001101,  // 0.8453295230865479
9'b000001110,  // 0.898597240447998
9'b000000100,  // 0.2548799514770508
9'b000001111,  // 0.9735668301582336
9'b000010010,  // 1.1261906623840332
9'b000000111,  // 0.44768181443214417
9'b111011010   // -2.3676068782806396
};
endpackage