// Width: 25
// NFRAC: 12
package dense_4_25_13;

localparam logic signed [24:0] weights [32][5] = '{ 
{25'b1111111111111111111001111, 25'b0000000000000010100001100, 25'b1111111111111101100111011, 25'b0000000000000000100001101, 25'b1111111111111111001001100}, 
{25'b1111111111111011100010011, 25'b1111111111111111100011110, 25'b0000000000000011101011101, 25'b1111111111111111111001101, 25'b0000000000000000001000100}, 
{25'b0000000000000010111110001, 25'b0000000000000001101100011, 25'b1111111111111111110001101, 25'b1111111111111100110000011, 25'b1111111111111110010100000}, 
{25'b1111111111111100111111101, 25'b1111111111111101000001000, 25'b1111111111111111000110110, 25'b0000000000000010011101100, 25'b0000000000000001111000010}, 
{25'b0000000000000000111110100, 25'b0000000000000001000001111, 25'b0000000000000001010000011, 25'b1111111111111111110110101, 25'b1111111111110111111001011}, 
{25'b0000000000000010100111011, 25'b1111111111111100110110000, 25'b0000000000000001011100111, 25'b1111111111111110101101011, 25'b1111111111111110101000110}, 
{25'b1111111111111100110010100, 25'b0000000000000000010010001, 25'b1111111111111111111111111, 25'b0000000000000001011001001, 25'b0000000000000000100011010}, 
{25'b1111111111111111111111000, 25'b0000000000000010010001101, 25'b1111111111111100110111010, 25'b0000000000000001010011010, 25'b0000000000000001000101101}, 
{25'b0000000000000001010011101, 25'b1111111111111110101001010, 25'b0000000000000000000000101, 25'b1111111111111100010011101, 25'b1111111111111110000000101}, 
{25'b1111111111111111111111111, 25'b1111111111111101110111101, 25'b0000000000000001011011000, 25'b0000000000000011011100001, 25'b0000000000000000000000000}, 
{25'b1111111111111110111101011, 25'b1111111111111110110101111, 25'b0000000000000000000000000, 25'b0000000000000100101001101, 25'b1111111111111101110110111}, 
{25'b0000000000000001010110101, 25'b0000000000000001110101010, 25'b1111111111111101010001111, 25'b1111111111111111110001111, 25'b0000000000000000111110010}, 
{25'b0000000000000000000000000, 25'b0000000000000001010101110, 25'b0000000000000000000100100, 25'b1111111111111110010101100, 25'b1111111111111011000001000}, 
{25'b0000000000000001011010110, 25'b0000000000000000100000101, 25'b0000000000000011010110110, 25'b1111111111111111011100001, 25'b1111111111111100100100111}, 
{25'b0000000000000000101110011, 25'b1111111111111111100111010, 25'b1111111111111101000111011, 25'b1111111111111111101111000, 25'b0000000000000100010010100}, 
{25'b1111111111111100001101010, 25'b1111111111111110000010111, 25'b1111111111111110001110000, 25'b0000000000000011001100001, 25'b0000000000000000010000011}, 
{25'b0000000000000010110001000, 25'b1111111111111110101000000, 25'b1111111111111110111010100, 25'b1111111111111110001100011, 25'b1111111111111111100001010}, 
{25'b0000000000000001100011110, 25'b1111111111111111101011010, 25'b1111111111111100101100111, 25'b1111111111111111110000010, 25'b0000000000000000100100001}, 
{25'b0000000000000010000100010, 25'b0000000000000000010101010, 25'b1111111111111110010000011, 25'b0000000000000000000000000, 25'b1111111111111100111111100}, 
{25'b0000000000000001110110011, 25'b1111111111111111010011101, 25'b1111111111111110010011000, 25'b0000000000000001101010000, 25'b0000000000000000110000101}, 
{25'b0000000000000000100010101, 25'b1111111111111111110000011, 25'b0000000000000010011000010, 25'b1111111111111100100011010, 25'b1111111111111111110101000}, 
{25'b0000000000000000000000000, 25'b0000000000000000111100010, 25'b0000000000000011111001001, 25'b1111111111111011110110101, 25'b1111111111111011000011110}, 
{25'b1111111111111111001101101, 25'b0000000000000000111000001, 25'b0000000000000001011010101, 25'b1111111111111101001001010, 25'b0000000000000100001011011}, 
{25'b1111111111111111111111110, 25'b0000000000000001010100011, 25'b0000000000000010010000101, 25'b0000000000000000010011011, 25'b1111111111111011011011000}, 
{25'b1111111111111110101001010, 25'b0000000000000010111010100, 25'b1111111111111110001101100, 25'b0000000000000000000010111, 25'b0000000000000011000110101}, 
{25'b0000000000000000001101011, 25'b0000000000000010001000000, 25'b0000000000000000001111001, 25'b1111111111111010000001000, 25'b0000000000000100011000101}, 
{25'b1111111111111100010100101, 25'b1111111111111110000011010, 25'b0000000000000001101101101, 25'b0000000000000001111101001, 25'b0000000000000001100111010}, 
{25'b0000000000000000000010000, 25'b0000000000000001111011011, 25'b1111111111111111101101010, 25'b1111111111111110110010111, 25'b0000000000000000010000001}, 
{25'b1111111111111111001010101, 25'b0000000000000001111110000, 25'b1111111111111011111110000, 25'b0000000000000001000111000, 25'b1111111111111110101110111}, 
{25'b1111111111111111110110100, 25'b0000000000000001001000010, 25'b1111111111111110101001100, 25'b1111111111111100110010111, 25'b0000000000000100101111111}, 
{25'b0000000000000011100101110, 25'b0000000000000000100011110, 25'b0000000000000010100110001, 25'b1111111111111011010010000, 25'b1111111111111101011110101}, 
{25'b1111111111111111100001101, 25'b1111111111111100111010010, 25'b0000000000000010111011010, 25'b0000000000000000100100010, 25'b0000000000000001000001010}
};

localparam logic signed [24:0] bias [5] = '{
25'b1111111111111111100000001,  // -0.06223141402006149
25'b1111111111111111011111111,  // -0.06270556896924973
25'b1111111111111111011100000,  // -0.07014333456754684
25'b0000000000000000101010000,  // 0.0820775106549263
25'b0000000000000001101110010   // 0.2155742198228836
};
endpackage