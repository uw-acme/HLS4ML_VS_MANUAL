//Width: 25
//Int: 9
package dense_1_gen;

localparam logic signed [24:0] weights [16][64] = '{
{25'b0000000000100000101001010, 25'b1111111110101100100100111, 25'b1111111111101000110111101, 25'b1111111111100011000000111, 25'b1111111111001100001010001, 25'b0000000000001110001000000, 25'b1111111101111011010000111, 25'b0000000000000000000001000, 25'b0000000000000111011011111, 25'b0000000000100001101111000, 25'b0000000000000000011000010, 25'b1111111111001100001101111, 25'b1111111111111111110111010, 25'b0000000000011010110000110, 25'b0000000000000100010010100, 25'b1111111111011110100000110, 25'b0000000000011101110011001, 25'b0000000000000111100000100, 25'b0000000000000000000000101, 25'b1111111111111111111110111, 25'b0000000000110000001111111, 25'b1111111111010101100100111, 25'b1111111111111101001011011, 25'b0000000000111100100000011, 25'b1111111111010110110110100, 25'b1111111110101000101000000, 25'b1111111111011100101111101, 25'b1111111111100111000000110, 25'b1111111111110010100111010, 25'b1111111111111111110001101, 25'b0000000000000100110101000, 25'b0000000000011111011010011, 25'b0000000000011001000011101, 25'b1111111111111110010100110, 25'b0000000000000000000001010, 25'b0000000000100111110111001, 25'b1111111111111101101100100, 25'b1111111111011111110110001, 25'b0000000000000011011111010, 25'b0000000000011000101001011, 25'b1111111111111110011101110, 25'b0000000000100011001110001, 25'b1111111111011101111001100, 25'b0000000001110110111000010, 25'b1111111111111111110111010, 25'b0000000000111001111011011, 25'b0000000000000000000000100, 25'b0000000000010111100110011, 25'b0000000000011001000110100, 25'b1111111111111100111111111, 25'b0000000000000000000000100, 25'b0000000000010100100010010, 25'b0000000000011011101001000, 25'b0000000000001001111101000, 25'b1111111111110001001111111, 25'b1111111111011000010001101, 25'b0000000001000100101010000, 25'b1111111111000000000011011, 25'b0000000000111011110111000, 25'b1111111111010010101001010, 25'b0000000001100101100001010, 25'b1111111111111111000011100, 25'b0000000000000001011101111, 25'b0000000000001010011000101},
{25'b0000000000000000010111001, 25'b1111111111010110111100001, 25'b1111111111101111000011000, 25'b1111111111011100001101111, 25'b1111111111010111010111110, 25'b0000000000001101101010000, 25'b1111111110011111011011101, 25'b1111111111111111101101101, 25'b1111111111100010111010001, 25'b0000000000010110000100010, 25'b0000000000000000110110001, 25'b1111111111110100111110001, 25'b0000000000011001001110111, 25'b0000000000000000000000100, 25'b1111111111111111111110111, 25'b0000000000011010100100111, 25'b1111111111111111001110111, 25'b0000000000000000000010110, 25'b1111111111101000101011101, 25'b1111111111011111111110011, 25'b0000000000111000100111111, 25'b1111111111110101101001001, 25'b0000000000000110001000110, 25'b0000000001011001011101010, 25'b0000000000100000111101110, 25'b1111111111100010100001011, 25'b1111111111100010011100011, 25'b1111111111111111111101010, 25'b1111111111110011000000111, 25'b1111111111001100000111111, 25'b1111111111111000010101101, 25'b0000000000111010001110100, 25'b0000000000100011101010010, 25'b0000000001000110011011000, 25'b0000000001010000100001001, 25'b0000000000000110011101101, 25'b1111111111110000110110001, 25'b1111111111001000011100100, 25'b0000000000000111010000001, 25'b0000000000011000001011011, 25'b0000000000000010111011111, 25'b0000000000011010011011010, 25'b1111111111100100110010011, 25'b0000000000100000010000010, 25'b0000000000010110000011111, 25'b0000000000000110011000010, 25'b1111111111010100011111011, 25'b0000000000001010001011011, 25'b0000000000100001010111110, 25'b0000000000000011110101100, 25'b0000000000000011001011100, 25'b0000000010010100001000010, 25'b1111111111110110011011111, 25'b1111111111110011011101001, 25'b1111111111111001000011001, 25'b1111111111111111000000011, 25'b0000000000100000111000110, 25'b1111111111010000101001101, 25'b0000000001111110000111111, 25'b0000000000000000100111011, 25'b0000000001000010101000110, 25'b0000000000011110101111110, 25'b0000000001101001010011101, 25'b0000000000010010000011011},
{25'b1111111111111111000001100, 25'b0000000000000000000000001, 25'b1111111111110101010110110, 25'b1111111111101001011110011, 25'b1111111111101000010111111, 25'b0000000000000101010110111, 25'b0000000010111101100011111, 25'b1111111111111111111111101, 25'b1111111101011101111100101, 25'b1111111111111111111111010, 25'b1111111111111111110001111, 25'b1111111111111101101101011, 25'b1111111111100010111001011, 25'b0000000000000000001010100, 25'b1111111111111110110011010, 25'b0000000000010101100001001, 25'b0000000001110011111001011, 25'b1111111111111111111111100, 25'b0000000000001001001111111, 25'b0000000000000000000010100, 25'b0000000000110100110000101, 25'b1111111110100011101011111, 25'b0000000001001001111010111, 25'b1111111110100100101001011, 25'b0000000001111001011010010, 25'b1111111111010011101010010, 25'b1111111111100000101010101, 25'b1111111110100100001001111, 25'b0000000010100011000001000, 25'b0000000000100011010011101, 25'b0000000000000001011101011, 25'b0000000001000010010001010, 25'b0000000010000010100111001, 25'b1111111101100111000011000, 25'b1111111111110011110001001, 25'b0000000000000100000101101, 25'b1111111111100010011011111, 25'b0000000001110010110100011, 25'b1111111111111010111101100, 25'b0000000000101000000100110, 25'b0000000000101010101000101, 25'b0000000000101111010100101, 25'b1111111111111111111111101, 25'b1111111111111111111110101, 25'b1111111111111101110010101, 25'b0000000000010100000111010, 25'b1111111111011100001100010, 25'b1111111111101010001101001, 25'b1111111111111101110001001, 25'b0000000000110010010110010, 25'b1111111111101001011110111, 25'b0000000000010011001110000, 25'b1111111111111111111100011, 25'b0000000000010001001011111, 25'b1111111111101001100010100, 25'b1111111111111111111111010, 25'b1111111111011000100010001, 25'b1111111110101010010011010, 25'b1111111111111111101111101, 25'b0000000000000000000000011, 25'b0000000011000101011111001, 25'b0000000000000001101010101, 25'b1111111111111111101010010, 25'b1111111111011000011001010},
{25'b1111111111000101010110110, 25'b1111111111010000110100100, 25'b1111111110100111010101101, 25'b0000000000100111011101001, 25'b1111111111010111100100011, 25'b1111111101010011101011101, 25'b1111111111110001010100100, 25'b1111111111011000100100100, 25'b0000000000011100101011100, 25'b1111111111111111111111111, 25'b0000000010100001111110010, 25'b1111111111110010011111110, 25'b1111111110011011110110011, 25'b0000000001001010001001001, 25'b0000000000000011001110010, 25'b1111111111111111110011110, 25'b1111111111000111001101000, 25'b1111111111111111111111101, 25'b0000000000000000000000110, 25'b1111111111100011000100000, 25'b1111111101101100101011101, 25'b1111111111110001101101100, 25'b1111111110100110100111101, 25'b0000000000011001011001110, 25'b1111111111001110011111001, 25'b1111111110001010001010001, 25'b0000000000101000000010011, 25'b0000000001011110010010010, 25'b0000000010100101110010110, 25'b1111111111000101001000000, 25'b1111111110110101011011000, 25'b0000000000001001011101000, 25'b0000000001000000000001100, 25'b1111111110010100010100000, 25'b1111111111010111110000001, 25'b0000000000000000000000000, 25'b1111111110100011000100100, 25'b0000000000011111000010101, 25'b1111111111000111100010011, 25'b0000000000001111010001111, 25'b0000000000111010101100110, 25'b0000000000010100000100010, 25'b0000000000000000000000000, 25'b0000000000000010100110100, 25'b0000000001000110101110011, 25'b1111111111100110011010001, 25'b1111111111111111111111001, 25'b1111111111010011111110100, 25'b1111111111111111111111000, 25'b1111111111110011100111101, 25'b1111111110110001001110100, 25'b0000000000001011000111000, 25'b1111111111111111111111011, 25'b0000000000011011111011001, 25'b0000000000101000010111110, 25'b0000000001010010110101011, 25'b1111111110000100001010000, 25'b1111111110001001000111011, 25'b1111111110100101110000000, 25'b0000000001101110111000001, 25'b0000000011011111111000111, 25'b1111111110001100110110011, 25'b1111111111111001000100110, 25'b0000000000110111100101101},
{25'b0000000000101011110011001, 25'b1111111110110000110101100, 25'b1111111111011110110011100, 25'b1111111111111111111111111, 25'b1111111111101100010010100, 25'b0000000000101011100011011, 25'b0000000000011000010000011, 25'b1111111111111111111110111, 25'b1111111110110011100010100, 25'b1111111111100001000100000, 25'b1111111111010000110011111, 25'b0000000000000110110001110, 25'b0000000000000000001010011, 25'b0000000000000000000000010, 25'b1111111111111010110100011, 25'b0000000000101101110010000, 25'b0000000000010001000110110, 25'b1111111111001101101101101, 25'b0000000000000011111011001, 25'b0000000000000001101110110, 25'b0000000000011010111001101, 25'b1111111111110000111001001, 25'b0000000000001001100001110, 25'b1111111111111101100011111, 25'b0000000010001000011011011, 25'b1111111111101000001001101, 25'b1111111111011100000000110, 25'b1111111111001100010101010, 25'b0000000000000000000000100, 25'b0000000000010101000101101, 25'b0000000000001110111000010, 25'b0000000000100011000001000, 25'b1111111111111110011010001, 25'b0000000000001001011111010, 25'b0000000000010000101110101, 25'b1111111111111111111111111, 25'b0000000000000000110010111, 25'b0000000001110000110101110, 25'b1111111111011011000001110, 25'b1111111111110110001100010, 25'b0000000000110111011101000, 25'b0000000000011111110110001, 25'b1111111111000001011010101, 25'b0000000000000000110000001, 25'b1111111101110111010000001, 25'b1111111111111111111111101, 25'b1111111111110000010100010, 25'b0000000000000001100001111, 25'b1111111111111111111110100, 25'b1111111111111101000000000, 25'b1111111111111111111111101, 25'b0000000000011000000100110, 25'b1111111111111111010110000, 25'b0000000000101000101011001, 25'b1111111111100111100010011, 25'b1111111110100001111001101, 25'b1111111111000100010011001, 25'b1111111110111110110011001, 25'b1111111110110001011011010, 25'b0000000001011111100110111, 25'b0000000010101111110101000, 25'b0000000001100101011111011, 25'b0000000000001111101100001, 25'b1111111111111111111110101},
{25'b1111111111000110111101111, 25'b1111111110101111010010001, 25'b0000000000000000000001000, 25'b0000000000100111010100110, 25'b0000000000100100100001000, 25'b1111111111100100110110111, 25'b0000000001001010100001011, 25'b1111111111111111111111001, 25'b0000000000011111001100000, 25'b1111111111111111111111101, 25'b1111111111111110110011011, 25'b1111111111110110101101010, 25'b1111111111101001011011000, 25'b0000000001001010000000011, 25'b1111111111110100100100111, 25'b0000000000000000000001101, 25'b1111111110110000000001010, 25'b1111111111010010101000111, 25'b0000000000000000000001000, 25'b1111111111111111111111000, 25'b1111111111111001111010011, 25'b1111111111010111110101010, 25'b1111111111010111001100110, 25'b0000000000111011100100110, 25'b1111111111010111010010101, 25'b1111111111111111111000110, 25'b0000000000100000110010001, 25'b1111111111110110101001100, 25'b1111111110001000100110110, 25'b1111111111111111111111011, 25'b1111111111110111011100010, 25'b1111111111111110101011111, 25'b1111111111111110100001001, 25'b0000000000000101001111001, 25'b0000000000010000111000100, 25'b0000000000101100010000001, 25'b0000000000000001101111100, 25'b1111111111110011011100101, 25'b1111111111011110011000111, 25'b1111111111111111110000101, 25'b1111111111101010010111010, 25'b1111111110111100111100110, 25'b0000000000110011001111101, 25'b0000000000000001011000001, 25'b0000000001001101001110111, 25'b0000000000000000000000001, 25'b1111111111111111111110111, 25'b0000000000001100001011000, 25'b1111111111001010010110100, 25'b0000000000011101111101001, 25'b0000000000000000000000001, 25'b1111111111110011000100001, 25'b1111111111010001101111110, 25'b0000000000110001011110011, 25'b1111111111111111111111111, 25'b0000000000101100011011001, 25'b0000000000011011101110101, 25'b0000000000011010000110011, 25'b1111111111111101100111010, 25'b1111111111111110111100011, 25'b1111111110011000100010101, 25'b1111111111101111110110000, 25'b1111111111111000101100011, 25'b1111111111111111111100110},
{25'b1111111111011011110011011, 25'b1111111111010101000110111, 25'b1111111111001000110000111, 25'b1111111111110111000110000, 25'b1111111111101110111100100, 25'b0000000000001101010110000, 25'b1111111110100110101000101, 25'b1111111111101100110010101, 25'b1111111111100011010010111, 25'b1111111111111111111110101, 25'b1111111111011011001101011, 25'b0000000000101100100010000, 25'b0000000000000100100011110, 25'b0000000000010001101000101, 25'b0000000000100111111100000, 25'b0000000000000000000010010, 25'b0000000001100110000010101, 25'b0000000000001011011100000, 25'b0000000000011111000101100, 25'b0000000000100010010111011, 25'b1111111111101011111100010, 25'b0000000000101110100000110, 25'b1111111111100000111100000, 25'b1111111110111111110000011, 25'b0000000000010110001100000, 25'b0000000001000010001001011, 25'b1111111111111111011101111, 25'b0000000000000110111001011, 25'b1111111110000110010010101, 25'b0000000000100100101011010, 25'b0000000000100010001100101, 25'b1111111111010000001110000, 25'b0000000000111100010110011, 25'b0000000001010101000101000, 25'b0000000000000000000000011, 25'b0000000000101011110100101, 25'b1111111111111111111111101, 25'b0000000000100100011000111, 25'b0000000000011001011111100, 25'b0000000000000000000000000, 25'b1111111111110000111010010, 25'b1111111111010001011101000, 25'b0000000000010010010111010, 25'b0000000000111101110111111, 25'b0000000001000010011100010, 25'b1111111111101010011110101, 25'b1111111111110101010100010, 25'b1111111111100111101100101, 25'b1111111111101110101100001, 25'b0000000000001111001001111, 25'b0000000000000000011010010, 25'b0000000000000100010111011, 25'b0000000000000000000000010, 25'b0000000000010111001110000, 25'b1111111111101001101010100, 25'b0000000001100010101011010, 25'b0000000000101101100100100, 25'b1111111111111100110101111, 25'b0000000000110001111101011, 25'b0000000000011011110010001, 25'b1111111100110000000000000, 25'b1111111110110110001111010, 25'b1111111111101001111101001, 25'b1111111111111110101110000},
{25'b0000000000000000101010001, 25'b0000000000011110100111111, 25'b1111111111111111111101010, 25'b1111111111111111111011110, 25'b1111111111010110110001000, 25'b1111111111111100000000100, 25'b1111111111011111000100000, 25'b0000000000000000000001000, 25'b0000000000000011100001111, 25'b0000000000110001110001011, 25'b0000000000000001110111110, 25'b1111111111001111101000001, 25'b1111111111110111111111111, 25'b0000000000000000000001011, 25'b1111111111111001010000001, 25'b1111111111000110011100110, 25'b1111111110010011011001111, 25'b1111111111111111111101110, 25'b1111111110110010101001101, 25'b1111111111000110111011100, 25'b1111111111001110001001001, 25'b0000000000101100011100010, 25'b0000000000000110000000100, 25'b1111111111101101110001010, 25'b1111111111001000000100011, 25'b0000000000010011111001001, 25'b0000000000000000000000010, 25'b0000000000111111111011000, 25'b0000000001100111001010101, 25'b1111111111111010110110101, 25'b0000000000000000000101111, 25'b0000000000011101100001000, 25'b1111111110101000101011100, 25'b1111111111010000100001110, 25'b0000000000000111000111000, 25'b0000000000001011110110101, 25'b1111111111011100000110000, 25'b0000000000011110101010010, 25'b0000000000010000111001111, 25'b1111111111101100011101000, 25'b1111111111001010010000111, 25'b1111111111111011010000110, 25'b0000000000000100001100110, 25'b1111111111101010101111010, 25'b0000000000000111001001001, 25'b0000000000011101010110111, 25'b1111111111110000101110001, 25'b0000000000000011000011110, 25'b0000000000000000000000011, 25'b1111111111100100000111111, 25'b1111111111001110010011111, 25'b0000000000110101010000000, 25'b0000000000010000001111111, 25'b1111111111101001001101000, 25'b0000000000010000111110000, 25'b1111111111111000000110100, 25'b1111111111000011010001011, 25'b1111111111101110111100011, 25'b1111111111111001010100001, 25'b1111111111110111000001100, 25'b0000000001101010010010110, 25'b0000000000011000011011111, 25'b1111111111111001110011001, 25'b1111111111111111111101011},
{25'b0000000000000001111000011, 25'b0000000001001011000111100, 25'b1111111110110101101011100, 25'b1111111111100010011011011, 25'b0000000000101001010011001, 25'b1111111111100101100111101, 25'b0000000010011011000010001, 25'b1111111111011011001011100, 25'b1111111111111111111110111, 25'b0000000000100101100010011, 25'b0000000000100000100010111, 25'b1111111111111111101011101, 25'b1111111111111001110110110, 25'b1111111111000010010010110, 25'b0000000000100100000001010, 25'b0000000000010100011100101, 25'b1111111111100111001100011, 25'b1111111111111111111111110, 25'b0000000000000000000000010, 25'b0000000000000000000010100, 25'b0000000000100001111101110, 25'b1111111111000101001010011, 25'b0000000000110010001100111, 25'b0000000001001110011100010, 25'b1111111111110100110101010, 25'b1111111111111111111101111, 25'b1111111111111101111010101, 25'b1111111111111111111110010, 25'b0000000001011110001111000, 25'b0000000000000000101000101, 25'b1111111111011101000001111, 25'b0000000000000000000000001, 25'b0000000000110001001011100, 25'b1111111110011000001100010, 25'b1111111110111010110010110, 25'b0000000000011001011100000, 25'b0000000000010001101110100, 25'b1111111110110110110110101, 25'b1111111111100111110010100, 25'b1111111111100100100101001, 25'b0000000000110011010101010, 25'b0000000000110010000010101, 25'b0000000000000000000000110, 25'b1111111111011101011100010, 25'b0000000000000000000110101, 25'b0000000000110010100111001, 25'b1111111111111000011101010, 25'b1111111111111111111110110, 25'b0000000000000001011110001, 25'b0000000000011111010111100, 25'b1111111111111000101001101, 25'b1111111111100111001110000, 25'b0000000000101100000011110, 25'b1111111111100100011110101, 25'b0000000000100011110011011, 25'b0000000001001010110101101, 25'b0000000000000101000111111, 25'b0000000000100001101111100, 25'b1111111111001100110001101, 25'b1111111111010001000010000, 25'b0000000001101010011110110, 25'b1111111111101111100001000, 25'b0000000000000101111000011, 25'b1111111111110100000010001},
{25'b0000000000000010000100110, 25'b1111111111000110000101110, 25'b0000000000101111001101111, 25'b1111111111011011101010011, 25'b1111111111111111101000000, 25'b0000000000011011000100101, 25'b1111111110110101100000101, 25'b0000000000011000100000011, 25'b0000000000111110110010000, 25'b0000000000010011101111010, 25'b0000000000101110011000011, 25'b0000000000101001010010001, 25'b1111111111011000111111111, 25'b1111111111110110010010100, 25'b1111111111111001011011000, 25'b0000000000000000001001110, 25'b1111111110000101001010011, 25'b0000000000101001010111011, 25'b1111111111111011010111110, 25'b0000000000000011111110110, 25'b1111111111010010111000001, 25'b0000000000001000111100100, 25'b0000000000010011100110001, 25'b1111111111111111111101000, 25'b1111111111000101000101100, 25'b1111111111111001111000110, 25'b1111111111110101100000011, 25'b0000000010011111101110110, 25'b1111111110101011001101000, 25'b0000000000001000100000011, 25'b0000000000001100011010110, 25'b1111111111111000100001011, 25'b1111111111100011101110001, 25'b0000000000001110111011000, 25'b1111111111110101111111010, 25'b1111111111101110110011001, 25'b1111111111101001001110000, 25'b1111111111100101000111010, 25'b1111111111111101001011000, 25'b1111111111011001111011100, 25'b0000000000101001001100010, 25'b0000000000001111110011000, 25'b0000000000111111100101110, 25'b0000000000001011001110101, 25'b0000000000000100101110001, 25'b1111111111011010110001001, 25'b0000000000000000000000001, 25'b1111111111111111111110101, 25'b1111111111111111111100010, 25'b0000000000011000110100000, 25'b0000000000010110101101101, 25'b0000000000100101101111101, 25'b1111111111111111001110010, 25'b1111111111011010011100101, 25'b0000000000000001001001111, 25'b0000000000000000000001000, 25'b0000000000101001010001100, 25'b1111111111100110010010010, 25'b1111111110111001100010100, 25'b0000000001000111110110001, 25'b1111111111011010011000110, 25'b0000000010010100111110000, 25'b1111111111111101011101110, 25'b1111111111010010101000000},
{25'b1111111110110110010000000, 25'b1111111111111111110000101, 25'b1111111111001011100100110, 25'b0000000000011101011111110, 25'b0000000000100001101101101, 25'b1111111111110010111010000, 25'b0000000001000010001011100, 25'b1111111111101010001100011, 25'b1111111111000010101001001, 25'b1111111111010001000010001, 25'b1111111111011111110110010, 25'b1111111111000011000101110, 25'b1111111111100010101100111, 25'b0000000000011001001101100, 25'b0000000000000000000000100, 25'b0000000000000000000010001, 25'b0000000001101011110110010, 25'b1111111111111010011110010, 25'b1111111111111111110111011, 25'b0000000000110100101000111, 25'b0000000000100101011111000, 25'b1111111110110101111011100, 25'b1111111111001111000011110, 25'b0000000000011000001100101, 25'b1111111111001000111000100, 25'b1111111111111101010100010, 25'b1111111111011110110001101, 25'b1111111111010101001110101, 25'b1111111111001000001111001, 25'b0000000000100110101011101, 25'b0000000000011101001010001, 25'b1111111111101100000010101, 25'b1111111111110110101100111, 25'b1111111110000011010101011, 25'b1111111111101001011000101, 25'b0000000000000110010101001, 25'b1111111111101111011010111, 25'b1111111111011010000011001, 25'b1111111111111111100010100, 25'b0000000000001111001110100, 25'b1111111111110000110000010, 25'b1111111111111111101010110, 25'b1111111111111011100001101, 25'b1111111110101010111111111, 25'b0000000000000000000110111, 25'b0000000000000000000000011, 25'b0000000000101011100010001, 25'b1111111111110000000101111, 25'b0000000000110110001110111, 25'b1111111111100111100111000, 25'b0000000000100100110111101, 25'b1111111111111111110100011, 25'b0000000000011100111010000, 25'b1111111111001101111010110, 25'b1111111111111111111111110, 25'b0000000001000001100010010, 25'b0000000000101000000010000, 25'b0000000000100101011001000, 25'b0000000000000011001111100, 25'b1111111111001100110100100, 25'b1111111111011001101110100, 25'b1111111110101000001011111, 25'b1111111111111111110000111, 25'b0000000000001101101101101},
{25'b0000000000100111011111011, 25'b0000000000000000010101000, 25'b0000000000010000110010000, 25'b1111111111111111111111111, 25'b0000000000010011101001000, 25'b1111111111101110110000001, 25'b0000000000011110000011100, 25'b0000000000000101011011110, 25'b0000000000010001011000101, 25'b0000000000101011100001100, 25'b1111111111011110010010000, 25'b1111111111111101010110000, 25'b1111111111111110111100011, 25'b1111111111111110111000010, 25'b1111111110101011100010101, 25'b1111111111011001111000101, 25'b0000000001010000101101101, 25'b1111111111111100011011010, 25'b1111111111111001010101001, 25'b0000000000000000000010001, 25'b1111111111001111010101111, 25'b0000000000000001001010101, 25'b0000000000100000000111101, 25'b0000000000000100110111110, 25'b0000000000000100101101001, 25'b0000000000101011010100010, 25'b0000000000000000000000010, 25'b0000000000000100110100011, 25'b0000000000000000000000000, 25'b1111111111111001111100001, 25'b1111111111100110010011100, 25'b1111111110101010110001010, 25'b0000000000100001110100011, 25'b0000000000101011111001101, 25'b1111111111111100010000001, 25'b1111111111100001111101111, 25'b0000000000000000000000001, 25'b1111111110101100001101100, 25'b1111111111111010001001001, 25'b1111111111111111100101111, 25'b0000000000011001000110000, 25'b1111111111101111010010111, 25'b1111111111111111111111001, 25'b0000000001101100011101110, 25'b0000000000111001011000011, 25'b1111111111111111001111100, 25'b1111111111111111111101011, 25'b1111111111111111111111001, 25'b1111111111100001001110000, 25'b0000000000010010110100101, 25'b0000000000010010011100100, 25'b0000000000010110010111000, 25'b0000000000010100001001001, 25'b0000000000110001101100101, 25'b0000000000101100110001010, 25'b0000000001010100011010100, 25'b1111111111101110000110110, 25'b0000000000110010010110011, 25'b0000000000010011100011001, 25'b1111111111010110010011101, 25'b0000000000001110001100000, 25'b1111111111001110010010001, 25'b1111111111000111101101110, 25'b1111111111000000001011011},
{25'b0000000000000000000010101, 25'b0000000000011101001111011, 25'b1111111111100111000110000, 25'b0000000000000000000000101, 25'b1111111111111001101110100, 25'b1111111111111011101000111, 25'b1111111110101011011101010, 25'b1111111111111111111111010, 25'b0000000000100000011100000, 25'b0000000000011111111110110, 25'b0000000000011110011011100, 25'b1111111111001101000010101, 25'b1111111111110100100101010, 25'b0000000000100100010110101, 25'b1111111111111111111101100, 25'b0000000000000000100111001, 25'b1111111110010100010011100, 25'b1111111111111111111101011, 25'b0000000000101111101011111, 25'b0000000000001001000001101, 25'b0000000000011110011110100, 25'b1111111111110001001111110, 25'b0000000000011111111101000, 25'b0000000000110011110101011, 25'b1111111111010010100001101, 25'b1111111111011100001100110, 25'b1111111111111111010110001, 25'b1111111111110101101010001, 25'b0000000000001000100110111, 25'b0000000000000000000001000, 25'b1111111111111111111111100, 25'b0000000000101000001110011, 25'b1111111110100000000001110, 25'b0000000000101110010000100, 25'b0000000001000000001011100, 25'b0000000000001110111010111, 25'b0000000000001110011001100, 25'b1111111111110010001011111, 25'b0000000000001110101111100, 25'b1111111111110010010101110, 25'b1111111111011111110110010, 25'b1111111111111001100011101, 25'b0000000000010101000011100, 25'b0000000001011001100001100, 25'b1111111110010011100001111, 25'b1111111111000110111100101, 25'b0000000000011000100101110, 25'b1111111111110011011110001, 25'b0000000000111001101011001, 25'b1111111111100001110001101, 25'b1111111111010101101000010, 25'b1111111111011100001000011, 25'b1111111111111111111111110, 25'b0000000000001111011001010, 25'b1111111111101011110111100, 25'b1111111110010100111010000, 25'b1111111111101101101100101, 25'b1111111111111110101100011, 25'b0000000000000101100100100, 25'b1111111110110001111000110, 25'b0000000010001111010111110, 25'b1111111110111010010101001, 25'b0000000001000101010101100, 25'b0000000000010011100111001},
{25'b0000000000001010000001001, 25'b1111111111100111011101010, 25'b0000000001010000011010011, 25'b1111111111011001010011101, 25'b1111111111000100101100001, 25'b0000000000001011100000011, 25'b0000000000100111100110111, 25'b0000000000100110011111000, 25'b1111111111101001010010011, 25'b1111111111101011011100101, 25'b0000000000000110101110010, 25'b0000000000011101010100110, 25'b0000000000011110000100011, 25'b0000000000000110011011001, 25'b1111111111100101110111100, 25'b0000000000010000011100000, 25'b0000000000111100010000011, 25'b1111111111111110100100101, 25'b1111111111011100001100111, 25'b0000000000000000000001011, 25'b0000000000001001100001110, 25'b0000000000000010100110010, 25'b1111111111011010011110110, 25'b0000000000001110011101001, 25'b0000000001100100101111101, 25'b0000000000000001010010000, 25'b0000000000010111000111101, 25'b1111111110011010011110101, 25'b1111111111110110101100101, 25'b0000000000000001001100001, 25'b1111111111100110111000111, 25'b1111111111011000000111100, 25'b0000000000111010101010011, 25'b1111111111111100100110010, 25'b1111111111111011001011010, 25'b1111111111011000111100101, 25'b0000000000010001101110011, 25'b0000000000100101011001001, 25'b1111111111111110110001100, 25'b1111111111111010011100001, 25'b1111111111101000000111100, 25'b0000000000011101001110000, 25'b0000000000000000000000101, 25'b1111111110101000001001100, 25'b0000000000100111110101101, 25'b0000000000110011000100110, 25'b1111111111111111111110001, 25'b0000000000000011010000111, 25'b1111111111001000011101101, 25'b1111111111110110011010011, 25'b1111111111111111111111110, 25'b1111111111010111010110100, 25'b0000000000000000000000011, 25'b1111111111101001111001100, 25'b0000000000000111010101101, 25'b1111111110010111011010000, 25'b1111111111111111111111111, 25'b1111111111111111111000111, 25'b0000000000100011001110010, 25'b0000000001001000000100001, 25'b1111111110100111000011110, 25'b0000000001000010100101100, 25'b0000000000000100110000000, 25'b1111111111110110011101001},
{25'b0000000000100100110101110, 25'b0000000010011110110000111, 25'b0000000000111111011011001, 25'b0000000000100100100000001, 25'b1111111111000010110111001, 25'b1111111111010111010111001, 25'b1111111010110011010001001, 25'b1111111111000101100001000, 25'b0000000000110011100101010, 25'b1111111111111111111111010, 25'b0000000000100101101001010, 25'b0000000001101110011111111, 25'b0000000000001000111001111, 25'b0000000000000000101101000, 25'b1111111111111101110101000, 25'b0000000000000000000001011, 25'b1111111111100111110000001, 25'b1111111111100110000100100, 25'b0000000000011101011101011, 25'b1111111110111111101111110, 25'b1111111110101010111000110, 25'b1111111111110010110111100, 25'b1111111110110101010000001, 25'b0000000000000011110001000, 25'b1111111011011100100110101, 25'b0000000001101000010111101, 25'b0000000001111110100111011, 25'b0000000001001101010000101, 25'b1111111100100000110110011, 25'b1111111111010111111101110, 25'b1111111110100111111100010, 25'b1111111110010100000001011, 25'b1111111010111100110010001, 25'b0000000001010110100101100, 25'b1111111111111010011001110, 25'b0000000000101000110011110, 25'b0000000000000011000010001, 25'b1111111101001000100101010, 25'b0000000000000000000010010, 25'b0000000000000000000000101, 25'b0000000000000100000101011, 25'b0000000010000010011110010, 25'b1111111111100101110000101, 25'b1111111110101101011101100, 25'b0000000001110010110111100, 25'b1111111111000111001100101, 25'b1111111111010110011110111, 25'b1111111111001101110000111, 25'b0000000000111101000111001, 25'b0000000001000100000000000, 25'b1111111111110111010011011, 25'b1111111111010011010100111, 25'b1111111111111111101110110, 25'b1111111111110001100111101, 25'b0000000000000000000000101, 25'b1111111111001111101110001, 25'b0000000001001101101000100, 25'b0000000010001010110010010, 25'b0000000001011011000101100, 25'b1111111110001011101010010, 25'b1111111000100110000000001, 25'b0000000001110001010101010, 25'b0000000000001011110101001, 25'b0000000000101000100100011},
{25'b1111111111100001000101001, 25'b0000000000101011001011001, 25'b0000000000101000101001101, 25'b1111111111111111110011000, 25'b1111111111010000011001011, 25'b1111111111110100100001011, 25'b1111111111001110111001010, 25'b1111111111111000111000001, 25'b0000000000010011000101011, 25'b1111111111110110011001000, 25'b1111111111111100000011000, 25'b1111111111111010111111010, 25'b1111111111111111111010011, 25'b1111111111101000100010011, 25'b1111111111111100100101100, 25'b1111111111110011001010001, 25'b0000000000101000000111111, 25'b1111111111111111111111110, 25'b1111111110101101111100101, 25'b0000000000111011100001101, 25'b0000000001001100001101101, 25'b0000000000110101000100111, 25'b1111111111010111011010111, 25'b1111111111101110011101111, 25'b1111111111010011101110001, 25'b1111111111011010111001100, 25'b0000000000011101000011101, 25'b0000000000011101111100100, 25'b0000000000011100111100011, 25'b0000000000101110000011110, 25'b0000000000000100011000100, 25'b0000000000110001011010110, 25'b1111111111111010101001001, 25'b0000000000000000100111101, 25'b0000000000100110111111101, 25'b0000000000010000110101110, 25'b1111111111110111100011010, 25'b1111111111111110110010011, 25'b0000000000000000000000111, 25'b1111111111011010100011100, 25'b1111111111100011011010110, 25'b1111111111110001111000010, 25'b1111111111010010000011000, 25'b0000000000111001100100101, 25'b0000000000000000000010010, 25'b1111111111111111010010101, 25'b1111111111110101011011001, 25'b1111111111101101000110110, 25'b1111111110011000111000111, 25'b1111111111111011000010001, 25'b1111111111100011010001100, 25'b1111111111101101110111001, 25'b1111111111110011001110000, 25'b0000000000100001110110101, 25'b0000000001010111010011011, 25'b0000000000010111111111110, 25'b1111111111111110010011001, 25'b1111111111010100000110101, 25'b1111111111111100001111001, 25'b0000000000000000000010110, 25'b0000000000101001101011110, 25'b1111111111111101010010110, 25'b0000000000000101110111110, 25'b0000000000000000000000000}
};
localparam logic signed [24:0] bias [64] = '{
25'b1111111111111011001110000,
25'b0000000000100011000001000,
25'b1111111111110000001001111,
25'b1111111111110111110000000,
25'b0000000000000110111110110,
25'b0000000000001110111100001,
25'b0000000000010001011101100,
25'b0000000000001001100101000,
25'b0000000000000101111110111,
25'b1111111111100110001101101,
25'b1111111111110011010100001,
25'b0000000000010011010101011,
25'b1111111111110010111010101,
25'b1111111111101101010010110,
25'b1111111111110100111100001,
25'b0000000000010101010001000,
25'b1111111111110101010010111,
25'b1111111111111000101000011,
25'b1111111111111011110111100,
25'b1111111111111100010111100,
25'b0000000000010000001000011,
25'b1111111111111011010000011,
25'b0000000000011000110000000,
25'b0000000000000010101110000,
25'b0000000000111111110100010,
25'b0000000000000010000001110,
25'b1111111111110101011000011,
25'b0000000000001110001001110,
25'b0000000000000001100000001,
25'b1111111111110010000111101,
25'b0000000000100011000111111,
25'b0000000000001011110001101,
25'b0000000000100011000110010,
25'b0000000000100010101001000,
25'b1111111111100000001110000,
25'b0000000000001010000000100,
25'b1111111111111111010000111,
25'b0000000000001101111000111,
25'b0000000000010001011001011,
25'b1111111111110000100001110,
25'b1111111111111000101111110,
25'b0000000000001011111010110,
25'b0000000000000111000000110,
25'b0000000000000011110010011,
25'b1111111111011000000011011,
25'b1111111111110101001010100,
25'b1111111111101010100001110,
25'b0000000000010010111001011,
25'b1111111111100001110001001,
25'b0000000000001000010111011,
25'b1111111111101111100011001,
25'b1111111111101110010101011,
25'b1111111111101100100110011,
25'b0000000000001010001101110,
25'b0000000000010111001110001,
25'b1111111111111001000101010,
25'b1111111111111110101101101,
25'b0000000000001000011101101,
25'b0000000000000110011110000,
25'b0000000000000011011100000,
25'b0000000000000100001101000,
25'b0000000000010011111010100,
25'b1111111111011011010110010,
25'b1111111111110100110001101
};
endpackage