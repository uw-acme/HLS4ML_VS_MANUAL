//Width: 25
//Int: 9
package dense_4_gen;

localparam logic signed [24:0] weights [32][5] = '{
{25'b1111111111111110011110110, 25'b0000000000101000011001101, 25'b1111111111011001110111000, 25'b0000000000001000011011010, 25'b1111111111110010011001100},
{25'b1111111110111000100111101, 25'b1111111111111000111101111, 25'b0000000000111010111010100, 25'b1111111111111110011011010, 25'b0000000000000010001001000},
{25'b0000000000101111100011111, 25'b0000000000011011000110100, 25'b1111111111111100011010111, 25'b1111111111001100000111010, 25'b1111111111100101000000111},
{25'b1111111111001111111011010, 25'b1111111111010000010001001, 25'b1111111111110001101100011, 25'b0000000000100111011001111, 25'b0000000000011110000101010},
{25'b0000000000001111101001000, 25'b0000000000010000011110001, 25'b0000000000010100000110111, 25'b1111111111111101101010000, 25'b1111111101111110010110010},
{25'b0000000000101001110111001, 25'b1111111111001101100001000, 25'b0000000000010111001110010, 25'b1111111111101011010111011, 25'b1111111111101010001100111},
{25'b1111111111001100101000100, 25'b0000000000000100100011101, 25'b1111111111111111111111111, 25'b0000000000010110010010101, 25'b0000000000001000110101100},
{25'b1111111111111111110000010, 25'b0000000000100100011010101, 25'b1111111111001101110110000, 25'b0000000000010100110100111, 25'b0000000000010001011011001},
{25'b0000000000010100111010000, 25'b1111111111101010010100100, 25'b0000000000000000001010101, 25'b1111111111000100111011110, 25'b1111111111100000001010110},
{25'b1111111111111111111110001, 25'b1111111111011101111010110, 25'b0000000000010110110001001, 25'b0000000000110111000010001, 25'b0000000000000000000000001},
{25'b1111111111101111010111000, 25'b1111111111101101011111111, 25'b0000000000000000000000001, 25'b0000000001001010011010111, 25'b1111111111011101101111100},
{25'b0000000000010101101011110, 25'b0000000000011101010101011, 25'b1111111111010100011110001, 25'b1111111111111100011110100, 25'b0000000000001111100101011},
{25'b0000000000000000000000101, 25'b0000000000010101011101010, 25'b0000000000000001001001010, 25'b1111111111100101011001101, 25'b1111111110110000010001101},
{25'b0000000000010110101100001, 25'b0000000000001000001010110, 25'b0000000000110101101101000, 25'b1111111111110111000010010, 25'b1111111111001001001111100},
{25'b0000000000001011100111110, 25'b1111111111111001110101101, 25'b1111111111010001110111001, 25'b1111111111111011110001110, 25'b0000000001000100101001101},
{25'b1111111111000011010100001, 25'b1111111111100000101110110, 25'b1111111111100011100001111, 25'b0000000000110011000011101, 25'b0000000000000100000110111},
{25'b0000000000101100010000111, 25'b1111111111101010000001000, 25'b1111111111101110101000011, 25'b1111111111100011001000000, 25'b1111111111111000010101010},
{25'b0000000000011000111101101, 25'b1111111111111010110100011, 25'b1111111111001011001110100, 25'b1111111111111100000101001, 25'b0000000000001001000011000},
{25'b0000000000100001000101101, 25'b0000000000000101010100101, 25'b1111111111100100000110001, 25'b0000000000000000000000001, 25'b1111111111001111111010000},
{25'b0000000000011101100111111, 25'b1111111111110100111011001, 25'b1111111111100100110000111, 25'b0000000000011010100001100, 25'b0000000000001100001011000},
{25'b0000000000001000101010111, 25'b1111111111111100000111111, 25'b0000000000100110000110000, 25'b1111111111001000110101101, 25'b1111111111111101010001101},
{25'b0000000000000000000000000, 25'b0000000000001111000101110, 25'b0000000000111110010010010, 25'b1111111110111101101010100, 25'b1111111110110000111100101},
{25'b1111111111110011011011111, 25'b0000000000001110000010110, 25'b0000000000010110101011010, 25'b1111111111010010010100100, 25'b0000000001000010110111001},
{25'b1111111111111111111100111, 25'b0000000000010101000110110, 25'b0000000000100100001011110, 25'b0000000000000100110111001, 25'b1111111110110110110001111},
{25'b1111111111101010010101001, 25'b0000000000101110101000100, 25'b1111111111100011011000010, 25'b0000000000000000101110111, 25'b0000000000110001101011110},
{25'b0000000000000011010111010, 25'b0000000000100010000000011, 25'b0000000000000011110010001, 25'b1111111110100000010000110, 25'b0000000001000110001011001},
{25'b1111111111000101001010100, 25'b1111111111100000110100111, 25'b0000000000011011011010001, 25'b0000000000011111010011001, 25'b0000000000011001110100111},
{25'b0000000000000000100001001, 25'b0000000000011110110110110, 25'b1111111111111011010100111, 25'b1111111111101100101111001, 25'b0000000000000100000011001},
{25'b1111111111110010101010010, 25'b0000000000011111100000101, 25'b1111111110111111100000001, 25'b0000000000010001110000110, 25'b1111111111101011101110111},
{25'b1111111111111101101001110, 25'b0000000000010010000100000, 25'b1111111111101010011001111, 25'b1111111111001100101111100, 25'b0000000001001011111110100},
{25'b0000000000111001011101100, 25'b0000000000001000111100110, 25'b0000000000101001100010011, 25'b1111111110110100100000011, 25'b1111111111010111101010100},
{25'b1111111111111000011011010, 25'b1111111111001110100100110, 25'b0000000000101110110100100, 25'b0000000000001001000100010, 25'b0000000000010000010100101}
};
localparam logic signed [24:0] bias [5] = '{
25'b1111111111111000000010010,
25'b1111111111110111111110011,
25'b1111111111110111000001011,
25'b0000000000001010100000011,
25'b0000000000011011100110000
};
endpackage