// Width: 10
// NFRAC: 5
package dense_2_10_5;

localparam logic signed [9:0] weights [64][32] = '{ 
{10'b0000001000, 10'b0000000000, 10'b1111111001, 10'b1111111111, 10'b0000001000, 10'b0000000000, 10'b1111111011, 10'b1111111111, 10'b1111110111, 10'b0000000010, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b1111111001, 10'b1111111110, 10'b1111110111, 10'b0000000000, 10'b1111111111, 10'b1111111001, 10'b1111111010, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b0000000011, 10'b0000001100, 10'b0000000101, 10'b1111111111, 10'b0000000001, 10'b1111110010, 10'b0000000000}, 
{10'b1111111100, 10'b1111111011, 10'b1111111011, 10'b1111111110, 10'b1111111111, 10'b0000000001, 10'b1111111000, 10'b0000000000, 10'b0000000000, 10'b1111111101, 10'b0000000100, 10'b1111111110, 10'b1111111110, 10'b1111111001, 10'b0000000000, 10'b1111111110, 10'b0000000000, 10'b1111111001, 10'b0000000101, 10'b0000000111, 10'b1111111110, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b1111111101, 10'b0000001000, 10'b0000000111, 10'b0000000000, 10'b0000000000, 10'b1111110000, 10'b0000000000, 10'b0000000000}, 
{10'b0000000010, 10'b1111111100, 10'b1111111011, 10'b1111111110, 10'b1111111101, 10'b1111111101, 10'b1111111010, 10'b0000000000, 10'b1111111011, 10'b0000000000, 10'b0000000000, 10'b1111111101, 10'b0000000010, 10'b1111111101, 10'b1111111111, 10'b1111111110, 10'b0000000000, 10'b0000000011, 10'b0000000001, 10'b0000000111, 10'b0000000001, 10'b1111111101, 10'b0000000000, 10'b0000000001, 10'b1111111111, 10'b0000000110, 10'b0000000100, 10'b0000000011, 10'b1111111111, 10'b1111111011, 10'b1111111111, 10'b0000000011}, 
{10'b0000000100, 10'b0000000000, 10'b0000000001, 10'b1111111111, 10'b1111101111, 10'b0000000000, 10'b0000000000, 10'b0000000111, 10'b0000000111, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b0000000110, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b1111111010, 10'b1111111110, 10'b0000000001, 10'b1111111101, 10'b1111111111, 10'b0000000000, 10'b1111111110, 10'b0000000010, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b1111111001, 10'b0000001001}, 
{10'b1111101010, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b1111111110, 10'b1111111011, 10'b0000000001, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b0000000110, 10'b0000000000, 10'b0000001010, 10'b1111111111, 10'b0000000110, 10'b1111110011, 10'b0000000000, 10'b1111111100, 10'b0000000101, 10'b0000001000, 10'b0000000000, 10'b0000000001, 10'b0000000101, 10'b0000000111, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b0000000111}, 
{10'b0000000001, 10'b1111111111, 10'b0000000100, 10'b1111101011, 10'b1111010011, 10'b1111110100, 10'b0000001011, 10'b1111101100, 10'b1111111111, 10'b1111101010, 10'b1111101111, 10'b1111110101, 10'b0000001011, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b1111111011, 10'b1111111111, 10'b1111110000, 10'b0000000000, 10'b0000000101, 10'b1111111111, 10'b0000000000, 10'b0000001000, 10'b0000000001, 10'b1111111111, 10'b1111111111, 10'b0000000110, 10'b1111111110, 10'b0000000110}, 
{10'b1111111110, 10'b1111111010, 10'b1111111000, 10'b1111111110, 10'b1111110110, 10'b0000000010, 10'b1111111010, 10'b1111111011, 10'b1111110010, 10'b0000000001, 10'b1111111111, 10'b1111111010, 10'b0000000011, 10'b1111111111, 10'b1111111110, 10'b1111101110, 10'b1111111111, 10'b0000000010, 10'b0000000110, 10'b1111111010, 10'b1111111011, 10'b1111111101, 10'b1111111111, 10'b0000000000, 10'b1111111110, 10'b1111101011, 10'b1111110111, 10'b1111111110, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b1111111111}, 
{10'b1111111011, 10'b1111111101, 10'b1111111101, 10'b1111111000, 10'b1111111100, 10'b1111111111, 10'b0000000011, 10'b1111111101, 10'b0000000110, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b0000000111, 10'b0000000000, 10'b1111111111, 10'b1111111101, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b0000000001, 10'b1111111010, 10'b0000000000, 10'b1111111111, 10'b1111111101, 10'b1111111111, 10'b0000000000, 10'b1111111111}, 
{10'b1111110000, 10'b1111111110, 10'b1111110011, 10'b0000000011, 10'b0000001111, 10'b1111111111, 10'b1111111111, 10'b0000000111, 10'b1111110001, 10'b1111111110, 10'b0000000000, 10'b1111111001, 10'b1111111111, 10'b0000000010, 10'b1111111001, 10'b0000011000, 10'b1111111111, 10'b0000000001, 10'b0000000110, 10'b0000000111, 10'b0000000000, 10'b1111110101, 10'b0000000000, 10'b0000001101, 10'b1111111010, 10'b0000010110, 10'b1111111011, 10'b1111111001, 10'b1111110000, 10'b1111110001, 10'b0000000000, 10'b0000000001}, 
{10'b0000000000, 10'b1111111111, 10'b1111111101, 10'b0000000000, 10'b0000001001, 10'b1111111111, 10'b1111111101, 10'b0000000010, 10'b0000000011, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b1111111100, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b0000000010, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b0000000001, 10'b1111111011, 10'b0000000010, 10'b0000000111, 10'b1111111111, 10'b0000000000, 10'b0000000001, 10'b0000000010}, 
{10'b0000000011, 10'b0000000000, 10'b1111111100, 10'b1111110111, 10'b1111100110, 10'b0000000100, 10'b0000000000, 10'b1111100101, 10'b0000000001, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b1111110011, 10'b1111111111, 10'b0000000111, 10'b0000000100, 10'b0000000110, 10'b1111110001, 10'b1111110100, 10'b0000000011, 10'b1111111110, 10'b1111111110, 10'b0000001011, 10'b1111111100, 10'b1111111111, 10'b1111111111, 10'b0000000110, 10'b1111111111, 10'b0000000000}, 
{10'b1111111001, 10'b1111110000, 10'b0000000000, 10'b1111111111, 10'b0000001010, 10'b1111110111, 10'b1111111000, 10'b0000000011, 10'b1111111111, 10'b0000000100, 10'b0000000010, 10'b1111111101, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b1111110111, 10'b0000000101, 10'b0000000000, 10'b0000001001, 10'b0000000010, 10'b0000000000, 10'b1111111110, 10'b0000000100, 10'b1111111101, 10'b1111110110, 10'b1111111111, 10'b0000000101, 10'b1111111111, 10'b0000000000, 10'b1111111100, 10'b0000000100, 10'b0000001000}, 
{10'b0000000000, 10'b0000000000, 10'b0000000111, 10'b0000000000, 10'b1111111110, 10'b0000000101, 10'b0000000010, 10'b1111111111, 10'b0000000000, 10'b1111111011, 10'b1111111110, 10'b1111111010, 10'b1111111111, 10'b0000000001, 10'b1111111101, 10'b0000011010, 10'b0000000000, 10'b1111111100, 10'b1111111001, 10'b1111111111, 10'b0000000110, 10'b0000000100, 10'b0000000000, 10'b1111111111, 10'b0000000111, 10'b0000001000, 10'b0000001111, 10'b0000000000, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b1111111101}, 
{10'b1111111011, 10'b0000000001, 10'b0000000001, 10'b1111111000, 10'b1111110111, 10'b0000001111, 10'b0000000001, 10'b0000000000, 10'b1111111010, 10'b1111111101, 10'b0000000100, 10'b0000000010, 10'b0000000000, 10'b1111111101, 10'b0000001001, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b1111111110, 10'b0000000010, 10'b0000000000, 10'b0000000011, 10'b1111111111, 10'b0000000000, 10'b0000010101, 10'b1111111110, 10'b1111111111, 10'b1111111111, 10'b1111111100, 10'b1111111110, 10'b0000000101}, 
{10'b0000000001, 10'b0000000010, 10'b0000001010, 10'b1111111110, 10'b0000000011, 10'b0000001011, 10'b0000000000, 10'b1111111111, 10'b0000000011, 10'b1111111100, 10'b1111111111, 10'b1111111100, 10'b0000000000, 10'b0000001100, 10'b1111111111, 10'b0000000000, 10'b0000000111, 10'b0000000000, 10'b0000000000, 10'b1111110101, 10'b1111111000, 10'b1111111110, 10'b1111111111, 10'b1111111011, 10'b1111111110, 10'b1111111101, 10'b1111111001, 10'b1111111001, 10'b0000000000, 10'b0000000011, 10'b1111110011, 10'b0000000000}, 
{10'b1111110110, 10'b0000000000, 10'b1111111111, 10'b1111111110, 10'b1111111111, 10'b0000000100, 10'b1111111101, 10'b0000001000, 10'b1111110100, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b1111111101, 10'b0000000010, 10'b0000000101, 10'b1111111111, 10'b1111110111, 10'b1111111110, 10'b0000000011, 10'b0000000010, 10'b0000000000, 10'b0000000000, 10'b0000000010, 10'b1111111000, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b1111111011}, 
{10'b1111110101, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b0000000011, 10'b0000000000, 10'b0000000001, 10'b0000000001, 10'b0000000010, 10'b0000000010, 10'b0000000101, 10'b0000000000, 10'b1111111100, 10'b0000000000, 10'b0000001100, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b0000000011, 10'b0000000100, 10'b0000000000, 10'b0000000001, 10'b1111111111, 10'b1111111110, 10'b0000000000, 10'b1111111101, 10'b1111111011, 10'b0000000110, 10'b1111111111, 10'b0000000001, 10'b1111111001}, 
{10'b0000000000, 10'b1111111111, 10'b0000000001, 10'b0000000000, 10'b0000011101, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b0000000011, 10'b1111111101, 10'b0000000000, 10'b0000000000, 10'b0000000000, 10'b0000000100, 10'b0000000000, 10'b1111111011, 10'b1111111111, 10'b1111111101, 10'b0000001010, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b0000000010, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b0000000001}, 
{10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b0000000001, 10'b1111111110, 10'b1111111100, 10'b1111111110, 10'b0000001000, 10'b0000000000, 10'b0000000011, 10'b1111111111, 10'b0000000010, 10'b1111111110, 10'b1111111010, 10'b1111111001, 10'b0000000000, 10'b1111111111, 10'b1111111110, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b0000000010, 10'b0000000001, 10'b1111111011, 10'b0000000011, 10'b1111111010, 10'b0000000000, 10'b0000000000, 10'b1111111010, 10'b0000000000, 10'b0000000001, 10'b1111111111}, 
{10'b1111111111, 10'b1111111100, 10'b0000000000, 10'b1111111110, 10'b0000000110, 10'b1111111111, 10'b1111111111, 10'b0000000011, 10'b1111110011, 10'b0000000000, 10'b1111111110, 10'b1111111111, 10'b0000001011, 10'b0000000111, 10'b1111111100, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b1111111011, 10'b1111111100, 10'b0000000100, 10'b0000000000, 10'b1111111011, 10'b0000000000, 10'b1111111101, 10'b1111111110, 10'b0000000100, 10'b0000000000, 10'b1111111000}, 
{10'b0000010100, 10'b0000001010, 10'b1111111000, 10'b0000000000, 10'b1111110100, 10'b0000000000, 10'b0000000111, 10'b0000000000, 10'b0000000111, 10'b1111111111, 10'b1111111011, 10'b1111111101, 10'b0000000100, 10'b0000000000, 10'b1111111100, 10'b0000000100, 10'b0000010001, 10'b1111111011, 10'b1111110110, 10'b0000000000, 10'b1111111111, 10'b1111111010, 10'b1111111111, 10'b1111111111, 10'b0000000010, 10'b1111110100, 10'b0000000010, 10'b1111111111, 10'b0000000000, 10'b0000000011, 10'b1111111111, 10'b0000000001}, 
{10'b1111111101, 10'b1111111001, 10'b1111111110, 10'b1111111010, 10'b1111111111, 10'b0000000001, 10'b0000000000, 10'b1111111111, 10'b0000000001, 10'b1111111111, 10'b0000000000, 10'b1111111001, 10'b0000000011, 10'b0000000010, 10'b1111111100, 10'b0000001110, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b0000001010, 10'b1111110000, 10'b1111111100, 10'b1111111110, 10'b1111111111, 10'b0000000110, 10'b1111111110, 10'b0000000000, 10'b0000001111, 10'b1111101111, 10'b1111110100, 10'b0000000000}, 
{10'b0000000000, 10'b1111111110, 10'b1111111111, 10'b0000000000, 10'b1111101000, 10'b1111101100, 10'b0000000000, 10'b1111111111, 10'b1111110111, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b1111111110, 10'b1111111110, 10'b1111111101, 10'b1111111011, 10'b0000001001, 10'b0000000000, 10'b0000000001, 10'b1111111111, 10'b1111111101, 10'b0000000000, 10'b1111111101, 10'b0000000111, 10'b1111101100, 10'b0000000111, 10'b1111111111, 10'b1111111111, 10'b0000000110, 10'b1111111111, 10'b0000000111}, 
{10'b1111111111, 10'b0000000000, 10'b1111111110, 10'b0000000010, 10'b0000000001, 10'b1111110101, 10'b0000000000, 10'b0000000010, 10'b0000010010, 10'b1111111111, 10'b0000000000, 10'b0000000001, 10'b0000001011, 10'b1111111110, 10'b0000000000, 10'b0000000011, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b1111110111, 10'b0000000001, 10'b0000000010, 10'b0000000000, 10'b1111111111, 10'b0000000110, 10'b0000000000, 10'b0000000100, 10'b1111110010, 10'b0000000011, 10'b0000001100, 10'b0000000000}, 
{10'b1111110100, 10'b0000000110, 10'b1111110111, 10'b0000000011, 10'b1111111100, 10'b0000000000, 10'b0000001111, 10'b1111111000, 10'b1111110110, 10'b0000000101, 10'b1111111000, 10'b1111111111, 10'b1111111111, 10'b0000001011, 10'b1111111111, 10'b1111110110, 10'b1111111111, 10'b0000001110, 10'b1111110000, 10'b1111111111, 10'b0000001010, 10'b1111110100, 10'b0000000001, 10'b1111111111, 10'b0000001000, 10'b1111101111, 10'b1111110100, 10'b1111111001, 10'b1111111111, 10'b0000000011, 10'b0000000000, 10'b0000000101}, 
{10'b1111111101, 10'b0000000001, 10'b1111111111, 10'b0000000100, 10'b1111111110, 10'b0000000111, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b0000010000, 10'b0000000000, 10'b0000000110, 10'b0000000000, 10'b1111111001, 10'b1111111101, 10'b1111111111, 10'b1111111111, 10'b0000000001, 10'b1111111111, 10'b1111111010, 10'b1111111111, 10'b0000001001, 10'b0000001001, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b1111111100}, 
{10'b1111111101, 10'b0000000000, 10'b0000001000, 10'b0000000000, 10'b0000000000, 10'b1111111100, 10'b0000000000, 10'b1111100100, 10'b0000000110, 10'b0000000000, 10'b0000000000, 10'b1111110100, 10'b0000000000, 10'b1111111011, 10'b1111111110, 10'b0000000000, 10'b0000000000, 10'b0000000000, 10'b0000000011, 10'b0000000000, 10'b1111111111, 10'b0000001010, 10'b0000001100, 10'b1111111000, 10'b1111111011, 10'b0000000111, 10'b1111110110, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b0000000101}, 
{10'b1111111100, 10'b1111111111, 10'b1111111000, 10'b1111111001, 10'b1111111111, 10'b1111111011, 10'b0000000000, 10'b0000000010, 10'b1111111000, 10'b1111111101, 10'b1111111110, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b1111111110, 10'b0000000011, 10'b0000000111, 10'b0000000100, 10'b1111111011, 10'b0000000001, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b1111111101, 10'b0000000010, 10'b1111111101, 10'b0000000001, 10'b1111111111, 10'b1111110110, 10'b1111111111, 10'b0000000111}, 
{10'b1111111111, 10'b1111111101, 10'b0000000010, 10'b0000001000, 10'b0000000010, 10'b0000000010, 10'b0000000001, 10'b1111111001, 10'b1111111001, 10'b0000000010, 10'b0000000000, 10'b0000000001, 10'b0000000000, 10'b0000000000, 10'b0000000110, 10'b0000000000, 10'b1111111110, 10'b0000000011, 10'b1111111111, 10'b1111111110, 10'b0000000011, 10'b1111111100, 10'b1111111111, 10'b0000000100, 10'b0000000000, 10'b1111111100, 10'b1111111001, 10'b1111111111, 10'b1111110111, 10'b0000000001, 10'b0000000011, 10'b0000000000}, 
{10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b1111111110, 10'b1111111011, 10'b1111111011, 10'b0000000010, 10'b0000000000, 10'b1111111010, 10'b0000000101, 10'b1111111111, 10'b1111111111, 10'b1111111100, 10'b0000000000, 10'b0000000000, 10'b1111111110, 10'b1111111111, 10'b1111111110, 10'b1111111101, 10'b0000000000, 10'b1111111011, 10'b0000000011, 10'b1111111001, 10'b0000000000, 10'b0000000001, 10'b0000000011, 10'b0000000000, 10'b0000000000, 10'b0000001001, 10'b0000000001, 10'b0000000000, 10'b0000000010}, 
{10'b1111111111, 10'b0000001000, 10'b1111111111, 10'b1111111110, 10'b1111111001, 10'b1111111101, 10'b0000001101, 10'b1111101001, 10'b1111110100, 10'b1111111001, 10'b1111111000, 10'b1111110111, 10'b1111111111, 10'b0000001111, 10'b1111111111, 10'b0000000000, 10'b1111111001, 10'b0000001110, 10'b1111110010, 10'b0000000000, 10'b1111111111, 10'b1111110101, 10'b0000000000, 10'b1111111111, 10'b0000000001, 10'b1111111110, 10'b1111111011, 10'b1111111111, 10'b0000000101, 10'b0000000000, 10'b1111111101, 10'b0000000000}, 
{10'b0000001011, 10'b1111111100, 10'b0000000100, 10'b1111111110, 10'b0000000010, 10'b1111111111, 10'b1111111111, 10'b1111111101, 10'b0000000000, 10'b0000000010, 10'b1111111111, 10'b1111111110, 10'b1111111111, 10'b0000000111, 10'b0000000000, 10'b0000000001, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b1111110110, 10'b1111111111, 10'b0000000001, 10'b1111111100, 10'b1111111011, 10'b1111111111, 10'b1111111111, 10'b0000010001, 10'b1111110110, 10'b1111111100}, 
{10'b1111111110, 10'b1111111100, 10'b1111111101, 10'b0000000001, 10'b0000000100, 10'b1111111011, 10'b1111111111, 10'b1111111000, 10'b0000000001, 10'b0000000100, 10'b1111111001, 10'b1111110111, 10'b0000000000, 10'b1111101010, 10'b1111111101, 10'b1111111100, 10'b1111111001, 10'b1111111111, 10'b0000000100, 10'b0000000000, 10'b1111111110, 10'b1111111110, 10'b0000000000, 10'b0000000000, 10'b1111111110, 10'b1111100111, 10'b1111101110, 10'b1111110111, 10'b0000000001, 10'b0000000110, 10'b1111111111, 10'b0000000111}, 
{10'b1111111101, 10'b1111111001, 10'b0000000101, 10'b0000000010, 10'b0000000001, 10'b1111111101, 10'b1111111110, 10'b0000000011, 10'b0000010001, 10'b1111111010, 10'b1111111111, 10'b1111111111, 10'b0000000011, 10'b1111111110, 10'b1111111111, 10'b1111111111, 10'b1111111100, 10'b1111111111, 10'b0000000000, 10'b0000000111, 10'b1111111011, 10'b1111111111, 10'b0000000100, 10'b1111111111, 10'b0000000000, 10'b0000010000, 10'b0000001010, 10'b0000000000, 10'b0000000000, 10'b1111110010, 10'b1111111101, 10'b1111111111}, 
{10'b0000000000, 10'b0000000001, 10'b1111111111, 10'b0000000000, 10'b0000000111, 10'b1111110000, 10'b0000000000, 10'b1111111100, 10'b0000000101, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b1111111100, 10'b0000001000, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b1111110101, 10'b0000000001, 10'b0000000101, 10'b1111111111, 10'b0000000011, 10'b1111111111, 10'b0000000010}, 
{10'b1111111001, 10'b0000000000, 10'b1111110000, 10'b0000000000, 10'b1111111110, 10'b1111111110, 10'b1111111111, 10'b1111111101, 10'b1111111110, 10'b1111111101, 10'b0000000001, 10'b0000000000, 10'b1111111010, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b0000000010, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b0000001000, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b0000001010, 10'b0000000110, 10'b0000000001, 10'b1111111100, 10'b1111111111, 10'b0000000010, 10'b0000000001}, 
{10'b0000000001, 10'b0000000001, 10'b1111111111, 10'b0000000000, 10'b1111110001, 10'b0000000001, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b1111111010, 10'b1111111111, 10'b0000000000, 10'b1111111010, 10'b0000000000, 10'b0000000000, 10'b0000000000, 10'b0000000000, 10'b1111110100, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b0000000100, 10'b1111111111, 10'b0000000000, 10'b0000001110, 10'b0000001010, 10'b0000000000, 10'b0000000000, 10'b1111111000, 10'b0000000000, 10'b1111111111}, 
{10'b0000000010, 10'b0000000001, 10'b0000001000, 10'b1111111000, 10'b0000000100, 10'b0000000011, 10'b0000000000, 10'b0000000110, 10'b0000000000, 10'b1111111111, 10'b0000000001, 10'b0000000000, 10'b1111111111, 10'b0000000011, 10'b1111111111, 10'b1111111110, 10'b0000000000, 10'b0000000001, 10'b1111111110, 10'b0000000011, 10'b0000000001, 10'b1111101101, 10'b1111111100, 10'b0000000010, 10'b1111111111, 10'b1111101111, 10'b1111111011, 10'b1111111111, 10'b1111111111, 10'b1111111110, 10'b0000000000, 10'b1111111110}, 
{10'b0000000000, 10'b1111111111, 10'b1111111101, 10'b1111111010, 10'b0000000001, 10'b0000000000, 10'b0000000011, 10'b1111111111, 10'b0000000111, 10'b1111111111, 10'b0000000000, 10'b1111110101, 10'b1111111111, 10'b0000000100, 10'b1111111111, 10'b1111110111, 10'b0000000000, 10'b1111111111, 10'b0000001000, 10'b1111111111, 10'b1111110010, 10'b1111111111, 10'b0000001000, 10'b1111111111, 10'b1111111111, 10'b0000000100, 10'b1111111100, 10'b0000000010, 10'b0000000000, 10'b1111111001, 10'b0000000000, 10'b0000000000}, 
{10'b1111111001, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b0000001111, 10'b1111111100, 10'b1111111111, 10'b1111111111, 10'b1111111110, 10'b1111111110, 10'b0000000010, 10'b0000000100, 10'b1111111110, 10'b0000000111, 10'b0000000000, 10'b1111111111, 10'b1111110110, 10'b1111111111, 10'b0000000000, 10'b1111111101, 10'b0000000000, 10'b0000000001, 10'b0000000000, 10'b1111111111, 10'b1111111110, 10'b1111111001, 10'b1111110110, 10'b0000000000, 10'b1111111100, 10'b0000000001, 10'b1111111111, 10'b0000000010}, 
{10'b1111110010, 10'b1111111010, 10'b1111111011, 10'b0000000000, 10'b0000010010, 10'b1111111000, 10'b0000000000, 10'b1111111110, 10'b1111110010, 10'b0000000100, 10'b1111111111, 10'b0000010010, 10'b0000000000, 10'b1111111110, 10'b1111111111, 10'b0000000001, 10'b1111111111, 10'b0000000000, 10'b1111111110, 10'b0000001111, 10'b0000000001, 10'b1111111110, 10'b0000000011, 10'b1111111111, 10'b1111111111, 10'b1111111100, 10'b1111111110, 10'b1111110001, 10'b1111111011, 10'b1111111111, 10'b1111111111, 10'b1111111110}, 
{10'b0000000111, 10'b1111100110, 10'b1111101000, 10'b1111111010, 10'b0000010101, 10'b1111111111, 10'b1111110100, 10'b0000001000, 10'b0000000001, 10'b0000000000, 10'b0000000110, 10'b1111110111, 10'b0000000000, 10'b0000000000, 10'b1111111110, 10'b0000000000, 10'b1111111100, 10'b1111100010, 10'b0000000101, 10'b0000001011, 10'b0000001000, 10'b0000000000, 10'b0000000000, 10'b1111110011, 10'b1111101011, 10'b1111111111, 10'b1111110110, 10'b1111110001, 10'b1111111001, 10'b1111100011, 10'b0000001101, 10'b0000001101}, 
{10'b0000000000, 10'b0000000000, 10'b0000000000, 10'b0000000000, 10'b0000001000, 10'b1111111010, 10'b0000000000, 10'b0000000010, 10'b1111110100, 10'b0000000001, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b0000000111, 10'b0000000001, 10'b0000000000, 10'b0000000001, 10'b0000001010, 10'b1111111001, 10'b0000000000, 10'b1111111010, 10'b1111111111, 10'b0000001010, 10'b0000000000, 10'b1111111111, 10'b1111101110, 10'b1111111111, 10'b1111111011, 10'b1111111110, 10'b0000000000, 10'b0000000100, 10'b0000000011}, 
{10'b1111111110, 10'b0000000100, 10'b1111110110, 10'b0000000000, 10'b0000000110, 10'b1111111110, 10'b1111111111, 10'b0000000101, 10'b0000000000, 10'b1111111111, 10'b1111111101, 10'b0000000000, 10'b0000000000, 10'b1111111110, 10'b1111111100, 10'b1111111101, 10'b1111111110, 10'b1111111101, 10'b1111111100, 10'b0000000000, 10'b1111111111, 10'b1111111110, 10'b1111111101, 10'b0000001100, 10'b0000000000, 10'b1111110100, 10'b1111111111, 10'b0000000011, 10'b0000000000, 10'b0000000000, 10'b0000001000, 10'b1111111111}, 
{10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b1111111011, 10'b1111100100, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b1111101100, 10'b0000000010, 10'b1111111100, 10'b1111111111, 10'b0000000000, 10'b1111110100, 10'b1111111110, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b0000000001, 10'b0000001011, 10'b1111111100, 10'b1111110110, 10'b0000000000, 10'b1111110111, 10'b1111111100, 10'b1111111000, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b1111110000, 10'b1111111110, 10'b0000000111}, 
{10'b0000000011, 10'b0000000111, 10'b1111111111, 10'b0000000101, 10'b1111111001, 10'b1111111100, 10'b0000000011, 10'b0000000010, 10'b1111111110, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b1111110101, 10'b1111111111, 10'b0000000100, 10'b1111111100, 10'b0000000001, 10'b1111111111, 10'b1111111111, 10'b0000000110, 10'b1111110101, 10'b0000001000, 10'b0000000001, 10'b0000000000, 10'b0000000110, 10'b0000000000, 10'b1111111110, 10'b1111110011, 10'b1111111100, 10'b1111111010, 10'b0000000101}, 
{10'b0000000000, 10'b0000000000, 10'b1111110100, 10'b1111111111, 10'b0000000110, 10'b1111111011, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b0000000000, 10'b1111111001, 10'b0000000011, 10'b0000000000, 10'b0000000000, 10'b0000000001, 10'b1111111111, 10'b1111111011, 10'b0000000000, 10'b0000000000, 10'b1111111110, 10'b1111111111, 10'b0000001001, 10'b1111111111, 10'b0000000000, 10'b1111110110, 10'b1111110101, 10'b0000000111, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b0000001001}, 
{10'b1111110101, 10'b1111111111, 10'b1111111001, 10'b0000000000, 10'b1111110100, 10'b0000000000, 10'b1111111111, 10'b1111111101, 10'b1111101110, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b1111111110, 10'b1111111011, 10'b1111111100, 10'b0000000010, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b0000001010, 10'b1111111111, 10'b0000000100, 10'b0000000010, 10'b1111111011, 10'b0000000110, 10'b1111111110, 10'b0000000000, 10'b1111111111, 10'b0000010010}, 
{10'b1111110101, 10'b0000000000, 10'b0000000001, 10'b1111111111, 10'b0000000111, 10'b1111110110, 10'b1111111111, 10'b0000001000, 10'b0000000101, 10'b0000000000, 10'b1111111111, 10'b1111111101, 10'b1111111101, 10'b1111111101, 10'b1111111110, 10'b0000000010, 10'b1111111111, 10'b0000000000, 10'b0000000100, 10'b0000000000, 10'b0000000000, 10'b0000000000, 10'b0000001000, 10'b0000000001, 10'b0000000000, 10'b1111111100, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b0000000010}, 
{10'b1111111111, 10'b0000000000, 10'b1111111001, 10'b1111111101, 10'b0000001001, 10'b1111111111, 10'b1111111101, 10'b0000000111, 10'b1111111110, 10'b0000001001, 10'b0000000010, 10'b1111111100, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b1111111101, 10'b1111110111, 10'b0000001000, 10'b0000000100, 10'b0000010100, 10'b0000000110, 10'b0000000111, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b0000000001, 10'b0000000010, 10'b1111110010, 10'b1111111111, 10'b1111111111, 10'b1111111111}, 
{10'b0000000000, 10'b1111111101, 10'b1111111100, 10'b0000000000, 10'b1111111000, 10'b0000000000, 10'b0000000110, 10'b0000000011, 10'b0000000001, 10'b1111111100, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b1111111110, 10'b0000000110, 10'b1111111111, 10'b1111111111, 10'b1111110110, 10'b0000000000, 10'b1111111001, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b0000000000, 10'b0000000100, 10'b1111111101, 10'b1111111111, 10'b1111110001, 10'b0000000010}, 
{10'b0000001110, 10'b1111111111, 10'b0000000010, 10'b1111111100, 10'b1111111101, 10'b0000000001, 10'b0000000101, 10'b0000000000, 10'b0000010000, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b0000000011, 10'b1111111111, 10'b0000000001, 10'b0000000011, 10'b1111111111, 10'b1111110001, 10'b1111111110, 10'b1111111111, 10'b0000000011, 10'b0000000000, 10'b1111111111, 10'b0000000011, 10'b0000000000, 10'b1111110111, 10'b1111111100, 10'b0000000100, 10'b1111111111, 10'b0000001000, 10'b1111111111, 10'b1111111010}, 
{10'b0000000000, 10'b0000000011, 10'b1111111111, 10'b1111111110, 10'b1111110100, 10'b1111111111, 10'b0000000001, 10'b1111111110, 10'b0000000101, 10'b1111111110, 10'b1111111111, 10'b1111111110, 10'b1111111111, 10'b1111111110, 10'b0000000000, 10'b0000001010, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b0000000001, 10'b0000000100, 10'b0000000000, 10'b0000000000, 10'b0000000001, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b0000000000, 10'b0000000011}, 
{10'b1111110110, 10'b0000000100, 10'b0000000000, 10'b1111111100, 10'b1111110011, 10'b1111111111, 10'b0000000010, 10'b1111110011, 10'b0000010000, 10'b0000000010, 10'b0000000000, 10'b0000000011, 10'b0000000001, 10'b0000000000, 10'b0000001101, 10'b1111111101, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b1111110010, 10'b0000000000, 10'b0000000100, 10'b0000000001, 10'b0000000001, 10'b1111101010, 10'b1111110101, 10'b1111111000, 10'b0000000000, 10'b1111111111, 10'b0000001010, 10'b1111111001}, 
{10'b1111111111, 10'b1111111001, 10'b1111111100, 10'b1111110010, 10'b1111110111, 10'b0000001010, 10'b0000001001, 10'b1111111010, 10'b0000000001, 10'b1111111110, 10'b1111111100, 10'b1111110111, 10'b0000000011, 10'b1111110110, 10'b0000000110, 10'b1111111111, 10'b0000001010, 10'b1111111111, 10'b1111111111, 10'b1111111011, 10'b1111111110, 10'b1111111101, 10'b1111110111, 10'b0000000010, 10'b1111111111, 10'b1111111111, 10'b1111111000, 10'b0000001010, 10'b0000001000, 10'b1111111101, 10'b1111101011, 10'b0000000100}, 
{10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b1111111100, 10'b0000000000, 10'b0000000000, 10'b0000000010, 10'b0000000000, 10'b0000000011, 10'b1111111111, 10'b0000000000, 10'b0000000011, 10'b0000000000, 10'b0000000000, 10'b1111111011, 10'b1111111100, 10'b0000000000, 10'b0000000101, 10'b0000000001, 10'b0000000100, 10'b1111111111, 10'b1111111010, 10'b1111111111, 10'b0000000010, 10'b1111111111, 10'b0000000001, 10'b1111111111, 10'b0000000010, 10'b0000000000, 10'b0000000010, 10'b1111110011, 10'b1111111111}, 
{10'b0000001001, 10'b1111111111, 10'b0000000100, 10'b1111110110, 10'b1111111001, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b1111111011, 10'b0000000000, 10'b0000000000, 10'b0000000000, 10'b0000000000, 10'b1111111011, 10'b0000000100, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b0000000011, 10'b1111111001, 10'b0000000011, 10'b0000000100, 10'b0000000100, 10'b1111111111, 10'b0000010001, 10'b1111111011, 10'b0000001011, 10'b1111111110, 10'b1111110100, 10'b1111111010, 10'b0000000100}, 
{10'b1111101110, 10'b1111111111, 10'b1111111011, 10'b1111111111, 10'b0000001000, 10'b1111111010, 10'b1111111110, 10'b0000000111, 10'b0000000011, 10'b1111111000, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b0000000100, 10'b1111111000, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b1111111001, 10'b1111111111, 10'b0000000000, 10'b1111110101, 10'b0000000010, 10'b0000010011, 10'b0000001011, 10'b1111111110, 10'b1111111010, 10'b1111110001, 10'b0000000000, 10'b1111111110}, 
{10'b0000000000, 10'b0000000110, 10'b0000000000, 10'b1111111011, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b0000000110, 10'b0000000110, 10'b1111111011, 10'b0000000100, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b1111111010, 10'b0000001000, 10'b1111111110, 10'b1111110101, 10'b0000000011, 10'b1111111111, 10'b1111111111, 10'b0000000011, 10'b1111111101, 10'b1111111111, 10'b1111111110, 10'b0000000010, 10'b1111111011, 10'b0000000100, 10'b1111110100, 10'b0000000010, 10'b1111111111, 10'b0000000101}, 
{10'b1111111110, 10'b0000000000, 10'b0000000010, 10'b0000000000, 10'b1111111110, 10'b1111111111, 10'b0000000011, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b0000000000, 10'b0000000000, 10'b1111111100, 10'b0000000000, 10'b0000000011, 10'b0000000001, 10'b0000000011, 10'b1111111111, 10'b1111111111, 10'b0000000100, 10'b0000000111, 10'b1111111100, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b1111110001, 10'b1111111111, 10'b1111111101, 10'b1111111111, 10'b0000010010, 10'b0000000000, 10'b1111111001}, 
{10'b1111111111, 10'b1111111100, 10'b1111111111, 10'b0000000000, 10'b0000000010, 10'b1111111111, 10'b0000000000, 10'b1111111111, 10'b0000000010, 10'b1111111111, 10'b0000000000, 10'b0000000001, 10'b0000001001, 10'b1111111100, 10'b0000000000, 10'b1111100100, 10'b1111111111, 10'b1111111110, 10'b0000000000, 10'b1111111110, 10'b0000000010, 10'b1111111000, 10'b0000000011, 10'b0000000011, 10'b1111111111, 10'b1111101001, 10'b1111111000, 10'b1111111111, 10'b1111111111, 10'b0000001100, 10'b1111111111, 10'b0000000100}, 
{10'b0000000001, 10'b0000000000, 10'b0000000101, 10'b1111111100, 10'b1111111101, 10'b0000000111, 10'b1111111010, 10'b0000000001, 10'b1111110110, 10'b0000000000, 10'b0000000000, 10'b1111111101, 10'b0000000000, 10'b0000000000, 10'b1111111001, 10'b0000001101, 10'b1111111000, 10'b1111111111, 10'b0000000011, 10'b1111111111, 10'b0000000010, 10'b1111110000, 10'b0000001010, 10'b1111111111, 10'b1111111100, 10'b0000001111, 10'b0000000100, 10'b1111111010, 10'b1111111011, 10'b1111101110, 10'b1111111111, 10'b0000000000}, 
{10'b1111111111, 10'b0000000000, 10'b1111111110, 10'b1111110111, 10'b1111111111, 10'b1111110011, 10'b0000000000, 10'b0000001001, 10'b0000000111, 10'b0000000000, 10'b0000000000, 10'b1111111100, 10'b0000001010, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b0000001101, 10'b0000000000, 10'b1111111110, 10'b1111111110, 10'b1111110101, 10'b0000000100, 10'b0000000000, 10'b0000000000, 10'b0000000001, 10'b1111111101, 10'b1111110001, 10'b0000001000, 10'b1111110001, 10'b0000000001, 10'b1111111101, 10'b0000000000}, 
{10'b0000000001, 10'b0000000101, 10'b0000000000, 10'b1111111111, 10'b1111110001, 10'b0000000000, 10'b1111111111, 10'b0000000111, 10'b0000001000, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b0000000000, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b0000000101, 10'b1111111100, 10'b1111110010, 10'b1111111110, 10'b1111111100, 10'b1111111100, 10'b1111111101, 10'b1111111111, 10'b1111111101, 10'b1111111111, 10'b1111111111, 10'b0000000100, 10'b1111111111, 10'b0000001110}
};

localparam logic signed [9:0] bias [32] = '{
10'b0000101111,  // 1.474280834197998
10'b0000010110,  // 0.6914801001548767
10'b0000101110,  // 1.4406442642211914
10'b0000101101,  // 1.408045768737793
10'b0000011111,  // 0.9864811301231384
10'b0000011011,  // 0.8636202812194824
10'b1111101100,  // -0.6153604388237
10'b0000001111,  // 0.4839226007461548
10'b0000001111,  // 0.4862793982028961
10'b0000001011,  // 0.37162142992019653
10'b0000001110,  // 0.45989668369293213
10'b0000101001,  // 1.2998151779174805
10'b1111011111,  // -1.016528844833374
10'b1111110100,  // -0.35249894857406616
10'b0000001110,  // 0.44582197070121765
10'b1111111100,  // -0.1119980737566948
10'b1111111101,  // -0.06717441976070404
10'b0000000000,  // 0.00487547367811203
10'b0000000110,  // 0.1946917623281479
10'b1111100111,  // -0.7796769738197327
10'b0000010111,  // 0.7287401556968689
10'b0000110110,  // 1.714877724647522
10'b1111001100,  // -1.5971007347106934
10'b0000000010,  // 0.07393483817577362
10'b0000001010,  // 0.3225609362125397
10'b0000011011,  // 0.8453295230865479
10'b0000011100,  // 0.898597240447998
10'b0000001000,  // 0.2548799514770508
10'b0000011111,  // 0.9735668301582336
10'b0000100100,  // 1.1261906623840332
10'b0000001110,  // 0.44768181443214417
10'b1110110100   // -2.3676068782806396
};
endpackage