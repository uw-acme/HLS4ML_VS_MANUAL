// Width: 28
// NFRAC: 14
package dense_3_28_14;

localparam logic signed [27:0] weights [32][32] = '{ 
{28'b1111111111111111110011011011, 28'b1111111111111110010000000100, 28'b1111111111111110011000001001, 28'b1111111111111111001111001111, 28'b0000000000000001010111110110, 28'b0000000000000000001011001111, 28'b1111111111111111111100101110, 28'b1111111111111111111111110010, 28'b1111111111111111111111111111, 28'b1111111111111111111111111101, 28'b0000000000000000100000010001, 28'b1111111111111101111001000111, 28'b1111111111111111110000101110, 28'b0000000000000011011000110110, 28'b1111111111111111000010001011, 28'b1111111111111100010001001110, 28'b1111111111111111110110101100, 28'b0000000000000000011100100001, 28'b0000000000000001101111010110, 28'b1111111111111110100110110101, 28'b1111111111111011101111001100, 28'b1111111111111111110100001111, 28'b0000000000000000001100100110, 28'b1111111111111110011000110000, 28'b0000000000000000000000000011, 28'b0000000000000100000011001111, 28'b1111111111111010001011001001, 28'b1111111111111111000111010000, 28'b1111111111111110011100100010, 28'b1111111111111111011001100101, 28'b0000000000000001101100010011, 28'b1111111111111111010111001101}, 
{28'b0000000000000010111111011010, 28'b0000000000000110111010111000, 28'b0000000000000001100110111011, 28'b1111111111111101010111101000, 28'b0000000000000000111110100010, 28'b1111111111111110111010000001, 28'b1111111111111111100100001110, 28'b0000000000000100010111000000, 28'b0000000000000000000001100001, 28'b1111111111111111111111111110, 28'b1111111111111111110111110111, 28'b1111111111111101101001011010, 28'b1111111111111111001100011100, 28'b0000000000000010001010010101, 28'b1111111111110111100100111010, 28'b1111111111111110000111010111, 28'b1111111111111111111111111111, 28'b1111111111111111111101111000, 28'b1111111111111111110010100001, 28'b1111111111111111010101111100, 28'b1111111111111110111101110110, 28'b1111111111111110111001100000, 28'b0000000000000000000100011010, 28'b1111111111111111111111100101, 28'b1111111111111111111110010110, 28'b1111111111111011101101100010, 28'b0000000000000000000011000000, 28'b0000000000000001111000100100, 28'b1111111111111111101111110011, 28'b1111111111111101001111011010, 28'b0000000000000000000000101100, 28'b0000000000000000001001101100}, 
{28'b1111111111111100000011110010, 28'b0000000000000000101111001001, 28'b0000000000000000000010101111, 28'b0000000000000001010010100111, 28'b1111111111111101011110101000, 28'b0000000000000000000000001000, 28'b0000000000000000000000011011, 28'b1111111111111100101001001011, 28'b0000000000000010001001001100, 28'b1111111111111110111100111011, 28'b1111111111111110111101100101, 28'b1111111111111010000011010110, 28'b1111111111111110110000011001, 28'b0000000000000010000010110011, 28'b0000000000000001000011100010, 28'b1111111111111111111111100100, 28'b1111111111111111100010101110, 28'b1111111111111111111001111100, 28'b1111111111111100101111011110, 28'b0000000000000000000000110011, 28'b0000000000000000011111111010, 28'b0000000000000000010001101010, 28'b0000000000000000110101100011, 28'b0000000000000011100001010011, 28'b0000000000000000001001101100, 28'b1111111111111100110110001111, 28'b0000000000000011000100011100, 28'b0000000000000000000000001011, 28'b0000000000000000101010011101, 28'b1111111111111111111010010111, 28'b0000000000000000000000001111, 28'b0000000000001001000100110101}, 
{28'b0000000000000011010110011100, 28'b1111111111111111111111111111, 28'b1111111111111111001110001111, 28'b0000000000000101001111000001, 28'b0000000000000100111010011000, 28'b0000000000000000000000000101, 28'b0000000000000000010010110111, 28'b0000000000000011010000010101, 28'b1111111111111110011010101001, 28'b1111111111111111111111111101, 28'b1111111111111100101101001111, 28'b0000000000000000011110101000, 28'b0000000000000001000100001110, 28'b1111111111111101000000101010, 28'b0000000000000000010111111100, 28'b1111111111111111010111000101, 28'b1111111111111111111111111101, 28'b1111111111111110100010110011, 28'b0000000000000000001001110110, 28'b0000000000000000001110001000, 28'b0000000000000000000100000100, 28'b1111111111111111101101010100, 28'b0000000000000100110001100101, 28'b0000000000000010101111100011, 28'b0000000000000010101000101000, 28'b0000000000000001111111000100, 28'b0000000000000010101110111001, 28'b0000000000000000000000000111, 28'b1111111111111111100001110010, 28'b0000000000000011100111111110, 28'b0000000000000001111111110001, 28'b1111111111111111010011000011}, 
{28'b0000000000000100000000001000, 28'b1111111111111111101000000101, 28'b1111111111111101001110100011, 28'b1111111111111001111111001101, 28'b0000000000000011110100011101, 28'b0000000000000000000000000100, 28'b1111111111111100101101111111, 28'b1111111111111101101111010011, 28'b1111111111111111101000001010, 28'b1111111111111001100001101011, 28'b1111111111110111001010010101, 28'b0000000000000011110010000001, 28'b0000000000000101010110011010, 28'b0000000000000100001011111100, 28'b1111111111111011011001100101, 28'b1111111111111001110011001101, 28'b0000000000000000000000000010, 28'b1111111111111110110111100110, 28'b0000000000000001100110110001, 28'b0000000000000001000111000001, 28'b1111111111111110011111100011, 28'b1111111111111111111100101111, 28'b0000000000000101110001011111, 28'b1111111111110101000000001000, 28'b0000000000000000101101000100, 28'b1111111111111010101110110100, 28'b0000000000000000100001100011, 28'b1111111111111110000000111101, 28'b1111111111111101100111001100, 28'b1111111111111111111111110101, 28'b0000000000000000100011110101, 28'b0000000000000100101001001110}, 
{28'b0000000000000000010110000111, 28'b1111111111111111101010110101, 28'b1111111111111101100010110011, 28'b1111111111111101111010101110, 28'b0000000000000010111110010100, 28'b0000000000000000000000000101, 28'b1111111111111101110000110000, 28'b1111111111111110111010010011, 28'b1111111111111100100100110010, 28'b1111111111111111011111001101, 28'b1111111111111111111111110000, 28'b0000000000000001010010000101, 28'b0000000000000000000000000000, 28'b0000000000000010110111001011, 28'b1111111111111011111101000010, 28'b1111111111111110111110101001, 28'b0000000000000000101101100110, 28'b1111111111111101101001111111, 28'b1111111111111110011010110111, 28'b1111111111111111111111111101, 28'b0000000000000000000110001111, 28'b0000000000000010011001011011, 28'b0000000000000011101111000111, 28'b1111111111111111111010100010, 28'b1111111111111111111111110010, 28'b0000000000000011001101001010, 28'b1111111111111011100110101001, 28'b1111111111111111111111111100, 28'b1111111111111110000110111001, 28'b1111111111111111101101001001, 28'b1111111111111111111110011000, 28'b0000000000000000000011010100}, 
{28'b0000000000000000100001010100, 28'b1111111111111101010101110011, 28'b0000000000000000110111011110, 28'b1111111111111111101100010011, 28'b1111111111111111111100001001, 28'b0000000000000001001101100001, 28'b1111111111111111001001101111, 28'b1111111111111010100101010101, 28'b1111111111111111111111111101, 28'b1111111111111110010101010100, 28'b1111111111111100010110001001, 28'b0000000000000011110001110001, 28'b0000000000000000000011101001, 28'b0000000000000101011110011001, 28'b0000000000000110101000010010, 28'b0000000000000000000001010101, 28'b1111111111111111111111111111, 28'b1111111111111101011110100100, 28'b1111111111111111100000010010, 28'b0000000000000010001011111101, 28'b1111111111111001111111111101, 28'b0000000000000001001111110111, 28'b0000000000000010100111000100, 28'b0000000000000000001001101111, 28'b0000000000000001001100110111, 28'b0000000000001001111100100100, 28'b1111111111111100110110001101, 28'b1111111111111111010001100110, 28'b1111111111111110011110110010, 28'b0000000000000011111001011000, 28'b1111111111111111100110110100, 28'b1111111111111110101001010010}, 
{28'b1111111111111011001110101101, 28'b0000000000000000001100001100, 28'b1111111111111010111101110111, 28'b0000000000000011011110110100, 28'b0000000000001000001110010100, 28'b0000000000000000111011011100, 28'b0000000000000000000001111101, 28'b0000000000000000011000001010, 28'b1111111111111111111111111111, 28'b0000000000000001000001100001, 28'b0000000000001010011010001001, 28'b1111111111111111111111110110, 28'b0000000000000011000011001011, 28'b0000000000000100111110111100, 28'b0000000000000110001001100001, 28'b0000000000001000011001101010, 28'b0000000000000000000000000001, 28'b1111111111111100001011001100, 28'b0000000000000010101100001011, 28'b1111111111111111111101001100, 28'b1111111111111010111001011011, 28'b1111111111111110001011110110, 28'b0000000000000000000110111001, 28'b1111111111111111010101100111, 28'b1111111111111011111111010100, 28'b0000000000001111000000010001, 28'b1111111111111110001111100100, 28'b0000000000000000000000000001, 28'b0000000000000000000000000001, 28'b0000000000000111000100000111, 28'b0000000000000000101101011001, 28'b0000000000000011001000100101}, 
{28'b0000000000000011011000001101, 28'b1111111111111111110110000011, 28'b0000000000000000000000001001, 28'b1111111111111111101001110100, 28'b0000000000000000101001110001, 28'b1111111111111111101100100000, 28'b1111111111111111111111110111, 28'b0000000000000001010000010101, 28'b0000000000000001101100001110, 28'b1111111111111101110011101110, 28'b0000000000000001000111101101, 28'b0000000000000001011111111100, 28'b0000000000000000000110000100, 28'b0000000000000010101010011000, 28'b1111111111111110001100110001, 28'b1111111111111001100111111101, 28'b0000000000000000000000000001, 28'b1111111111111111111000110110, 28'b1111111111111111110010010101, 28'b1111111111111100000000101111, 28'b1111111111111111111111011011, 28'b0000000000000000000000000011, 28'b1111111111111110011000001100, 28'b1111111111111111111000110001, 28'b1111111111111111001111010111, 28'b0000000000000001001111110000, 28'b0000000000000010111111010101, 28'b1111111111111111000010110100, 28'b1111111111111111100110110110, 28'b1111111111111111101011011001, 28'b0000000000000000001101110101, 28'b1111111111111100110111000101}, 
{28'b1111111111111110100101000010, 28'b0000000000000011000100110100, 28'b0000000000000000000000000011, 28'b0000000000000000000000000001, 28'b0000000000000110010101101010, 28'b0000000000000010100100111110, 28'b1111111111111111111111111111, 28'b1111111111111011100011110011, 28'b0000000000000000111100010110, 28'b1111111111111010011010110101, 28'b1111111111110100110001100111, 28'b1111111111111111111111111101, 28'b0000000000000000000000001010, 28'b0000000000000011011011101000, 28'b0000000000000000111000110100, 28'b0000000000000000000000000010, 28'b1111111111111101010111110100, 28'b0000000000000000000000001011, 28'b0000000000000000000011011100, 28'b0000000000000000011111000010, 28'b0000000000000001111100110101, 28'b1111111111111111110010111110, 28'b1111111111111101000111100101, 28'b0000000000000000000100001101, 28'b1111111111111111111010001101, 28'b0000000000001000101001101100, 28'b0000000000000010100111001110, 28'b1111111111111111111111110011, 28'b1111111111111111011011101110, 28'b0000000000000101010110001011, 28'b1111111111111111101011100111, 28'b1111111111111111010011001011}, 
{28'b1111111111111011110100001111, 28'b0000000000000001011001101111, 28'b1111111111111111101110001111, 28'b1111111111111111111111111101, 28'b1111111111111110000001111100, 28'b1111111111111100111110101001, 28'b0000000000000000011000100110, 28'b0000000000000001001001110101, 28'b1111111111111111111111111111, 28'b1111111111111110101000010111, 28'b1111111111111011011010110101, 28'b0000000000000001100110110100, 28'b0000000000000010011011101110, 28'b0000000000000000000000000001, 28'b0000000000000110101101100011, 28'b1111111111111011100000011000, 28'b0000000000000000110101001110, 28'b1111111111111100110111110011, 28'b0000000000000010010000011000, 28'b1111111111111111111111111000, 28'b1111111111111111101100010001, 28'b0000000000000000100011111110, 28'b0000000000000000111110110100, 28'b0000000000000000000000000100, 28'b1111111111111100000011001110, 28'b0000000000000000001111111011, 28'b1111111111111011100001111001, 28'b1111111111111111101011101001, 28'b1111111111111111111111111000, 28'b0000000000000101011001111111, 28'b1111111111111110011110101011, 28'b0000000000000000000000001001}, 
{28'b1111111111111111111111111101, 28'b0000000000000000111010110011, 28'b0000000000000000000000001000, 28'b0000000000000011001000010101, 28'b1111111111111111000100000011, 28'b1111111111111111101001111100, 28'b0000000000000000011101111110, 28'b1111111111111111111101000001, 28'b1111111111111111101000010011, 28'b0000000000000101001000000000, 28'b0000000000000101100101111100, 28'b0000000000000000000000010110, 28'b1111111111111101010101101111, 28'b1111111111111010011000011100, 28'b1111111111111111100110000010, 28'b0000000000000000000000000101, 28'b0000000000000000000000000101, 28'b1111111111111111011111011000, 28'b1111111111111100001100000010, 28'b0000000000000011000011110001, 28'b0000000000000000000001000100, 28'b0000000000000010111101111100, 28'b1111111111111111111111111000, 28'b0000000000000100011111111110, 28'b0000000000000000111111010110, 28'b0000000000000010011100110110, 28'b0000000000000011101001001111, 28'b1111111111111111100101100001, 28'b1111111111111100110111100101, 28'b1111111111111100011110011001, 28'b1111111111111111111101011010, 28'b1111111111111010101001100001}, 
{28'b1111111111111110001100000111, 28'b1111111111111111111111111110, 28'b0000000000000000111101000100, 28'b1111111111111100101001100000, 28'b0000000000000000101100000110, 28'b1111111111111111111111111100, 28'b1111111111111110010000110011, 28'b1111111111111111111011000100, 28'b1111111111111110111111110011, 28'b0000000000000000010011000001, 28'b0000000000000000100111111010, 28'b1111111111111111011011011011, 28'b0000000000000000001000011100, 28'b0000000000000001100000000100, 28'b1111111111111010111111111110, 28'b1111111111111110000010101111, 28'b0000000000000001110100110100, 28'b1111111111111110100101011011, 28'b0000000000000000000000000010, 28'b1111111111111111110011001001, 28'b0000000000000001100010110011, 28'b0000000000000000000100000110, 28'b1111111111111111110000000100, 28'b0000000000000000010101110000, 28'b0000000000000010001001111101, 28'b1111111111111111001010110011, 28'b0000000000000000000000000110, 28'b1111111111111100011000101110, 28'b1111111111111110011011110010, 28'b1111111111111111111100011010, 28'b0000000000000001011000110001, 28'b0000000000000000000000001011}, 
{28'b1111111111111011110101111000, 28'b0000000000000011010111001110, 28'b1111111111111111111111111110, 28'b1111111111111111111100100101, 28'b1111111111111111111011000100, 28'b0000000000000001011001110001, 28'b1111111111111111111111111000, 28'b0000000000000110001011010011, 28'b1111111111111111111000011011, 28'b1111111111111111111111111110, 28'b0000000000000001101001011000, 28'b0000000000000000010100111111, 28'b0000000000000000000011010101, 28'b0000000000000000000000000111, 28'b0000000000000000111110010110, 28'b0000000000000010101001000011, 28'b0000000000000001011011001110, 28'b0000000000000001010101010111, 28'b1111111111111111111011101000, 28'b0000000000000010011101010011, 28'b0000000000000000110011100010, 28'b0000000000000000010100101111, 28'b1111111111111111111011100110, 28'b0000000000000010000010000010, 28'b1111111111111111001101000000, 28'b1111111111111101010010011111, 28'b1111111111111111010000101101, 28'b1111111111111111111111111110, 28'b0000000000000000110100000001, 28'b0000000000000000001111001101, 28'b0000000000000001100100000010, 28'b0000000000000011110101010100}, 
{28'b1111111111111111110110011100, 28'b1111111111111100111000101011, 28'b0000000000000000011010011100, 28'b1111111111111111111111100000, 28'b0000000000000111010101000010, 28'b1111111111111110010101110101, 28'b1111111111111011011011010110, 28'b0000000000000000000000000110, 28'b0000000000000000000000000011, 28'b1111111111111111110010110010, 28'b0000000000000000011000110011, 28'b0000000000000011011111100111, 28'b0000000000000010100100110101, 28'b0000000000000000000101011101, 28'b0000000000000000010001000100, 28'b1111111111111110100110100010, 28'b0000000000000000010001000100, 28'b1111111111111111101100100100, 28'b0000000000000000000000000011, 28'b0000000000000000100110100110, 28'b1111111111111111101100110101, 28'b0000000000000000001001110011, 28'b0000000000000010001000010100, 28'b0000000000000000010010111000, 28'b1111111111111111111001110101, 28'b1111111111111100101100101100, 28'b0000000000000001101000000010, 28'b1111111111111111111111111101, 28'b1111111111111111111111110100, 28'b1111111111111111001001100100, 28'b1111111111111111110101000001, 28'b1111111111111111011111111101}, 
{28'b0000000000000000000011101000, 28'b1111111111111111011111100110, 28'b1111111111111110111111011100, 28'b1111111111111110010000000000, 28'b1111111111111011101000001001, 28'b0000000000000100111000000010, 28'b0000000000000000000000000111, 28'b0000000000000001010110011111, 28'b0000000000000010010010111100, 28'b0000000000000000000110100100, 28'b1111111111111111101110101011, 28'b0000000000000011110011100011, 28'b0000000000000001110010100111, 28'b1111111111111101000100110101, 28'b1111111111111110101100111000, 28'b1111111111111111101010111011, 28'b1111111111111100110100000000, 28'b1111111111111111110111000111, 28'b0000000000000000000000000110, 28'b1111111111111111111101101010, 28'b0000000000000001001111110111, 28'b1111111111111110111001111111, 28'b0000000000000000000000000001, 28'b0000000000000000100111011010, 28'b1111111111111111111111111101, 28'b1111111111111101010001000011, 28'b0000000000000001010000001111, 28'b0000000000000000000000001101, 28'b0000000000000000010110110111, 28'b0000000000000000000101100111, 28'b1111111111111101011110001011, 28'b0000000000000000001010101000}, 
{28'b1111111111111110011011100111, 28'b1111111111111110101111011011, 28'b0000000000000000100111001000, 28'b1111111111111111000000011101, 28'b1111111111111111010010000000, 28'b0000000000000000111011011111, 28'b1111111111111111111101011000, 28'b0000000000000000010001111000, 28'b0000000000000001000011000100, 28'b1111111111111111111111110100, 28'b0000000000000000111111010111, 28'b1111111111111110111110110101, 28'b1111111111111111111011000010, 28'b1111111111111111111111111010, 28'b0000000000000000110100111101, 28'b1111111111111111111111111101, 28'b0000000000000011111010000111, 28'b1111111111111111110111000111, 28'b0000000000000001111111000000, 28'b1111111111111110101001000101, 28'b0000000000000001010001000001, 28'b0000000000000000100000001011, 28'b0000000000000000101011001101, 28'b0000000000000000010010100100, 28'b1111111111111111010110010100, 28'b1111111111111101110001010000, 28'b1111111111111101111011010110, 28'b0000000000000000110111010000, 28'b1111111111111111010101001001, 28'b0000000000000000000000010010, 28'b1111111111111111110001111110, 28'b0000000000000001110110110101}, 
{28'b1111111111111111111111111101, 28'b1111111111111100110000101110, 28'b1111111111111100110100111110, 28'b1111111111111111111111111100, 28'b0000000000000101000011001111, 28'b1111111111111111010001100010, 28'b0000000000000000000000000101, 28'b0000000000000011110111011100, 28'b1111111111111110110100011111, 28'b0000000000000000000000000010, 28'b1111111111111100101010001000, 28'b1111111111111100000101000010, 28'b0000000000000011100101100001, 28'b0000000000000001001101011000, 28'b1111111111111111000001111001, 28'b1111111111111101110011110110, 28'b0000000000000001011000010001, 28'b0000000000000000000000001110, 28'b1111111111111110000110010010, 28'b0000000000000000001101100110, 28'b0000000000000000100011100110, 28'b1111111111111111010010101111, 28'b0000000000000010010001011010, 28'b1111111111111000001010011001, 28'b0000000000000000010100111111, 28'b0000000000000001111010011001, 28'b1111111111111111101010111011, 28'b0000000000000000000111101000, 28'b1111111111111110001000100100, 28'b1111111111111111111111111011, 28'b1111111111111110011001000000, 28'b1111111111111111110011101010}, 
{28'b0000000000000001101100110110, 28'b0000000000000010110000101110, 28'b0000000000000100011001111111, 28'b1111111111111110010111010010, 28'b0000000000000011010101000010, 28'b0000000000000010011100110101, 28'b0000000000000000000000010000, 28'b0000000000000011101001001100, 28'b0000000000000010110110110111, 28'b1111111111111111001001010011, 28'b0000000000000101100111001111, 28'b1111111111111101001101001101, 28'b0000000000000100111110001000, 28'b0000000000000011100100100011, 28'b1111111111110111011010101000, 28'b1111111111111111111111100000, 28'b0000000000000000000000000010, 28'b0000000000000000000010111100, 28'b0000000000000010000101000101, 28'b1111111111111011111110010111, 28'b0000000000000001110001011111, 28'b1111111111111110010011011111, 28'b1111111111111100000100111111, 28'b1111111111111110101111101100, 28'b0000000000000010101000101000, 28'b1111111111111010101110001100, 28'b1111111111111101010111001010, 28'b1111111111111111101010111010, 28'b1111111111111111111111111011, 28'b1111111111111011011111000101, 28'b0000000000000011001010011111, 28'b0000000000000000000000001100}, 
{28'b1111111111111111100110110000, 28'b0000000000000000000000010111, 28'b1111111111111111111111111110, 28'b1111111111111111111111111111, 28'b1111111111111101001100001101, 28'b0000000000000000000100101101, 28'b0000000000000000000100001110, 28'b1111111111111111111000010011, 28'b1111111111111111110011100111, 28'b1111111111111111101000011101, 28'b0000000000000001000111001010, 28'b1111111111111111111111100111, 28'b0000000000000000101010011101, 28'b1111111111111101010000110011, 28'b0000000000000000110110101111, 28'b1111111111111111111111101000, 28'b0000000000000001001000000011, 28'b0000000000000011100101001101, 28'b1111111111111101001011011010, 28'b0000000000000000011010100100, 28'b1111111111111111001101010001, 28'b0000000000000001000001110111, 28'b0000000000000001100001010110, 28'b1111111111111111010100010110, 28'b1111111111111101111111011000, 28'b0000000000000000001010100010, 28'b0000000000000110101000100110, 28'b1111111111111111110011100110, 28'b1111111111111111111000001011, 28'b0000000000000010100110000011, 28'b0000000000000000000000000110, 28'b0000000000000110111001010110}, 
{28'b1111111111111011110100111100, 28'b0000000000000000010010100000, 28'b1111111111111110010001001111, 28'b0000000000000011000100000011, 28'b0000000000000000111000001011, 28'b1111111111111111101111110100, 28'b1111111111111111111111111110, 28'b1111111111111111111111111111, 28'b1111111111111101100100110011, 28'b1111111111111111101111000111, 28'b0000000000000000000000000100, 28'b1111111111111011100011101100, 28'b0000000000000000000110011010, 28'b1111111111111111101011101001, 28'b1111111111111111111110101111, 28'b1111111111111111111111111001, 28'b1111111111111111000100010001, 28'b0000000000000000000010110010, 28'b0000000000000000000001100111, 28'b0000000000000001010001001111, 28'b0000000000000000001000111110, 28'b0000000000000000000000000001, 28'b0000000000000000000000000100, 28'b1111111111111111111011110110, 28'b0000000000000000000000001001, 28'b0000000000000000001001011000, 28'b0000000000000100101001101001, 28'b1111111111111111111111111110, 28'b1111111111111111111111111010, 28'b1111111111111111101011001001, 28'b0000000000000001011001101000, 28'b1111111111111111110010111101}, 
{28'b1111111111111111111111001100, 28'b1111111111111110110010100000, 28'b0000000000000001101000100110, 28'b0000000000000000010100011101, 28'b1111111111111101000001101011, 28'b0000000000000000000000010011, 28'b0000000000000010010010011010, 28'b1111111111111111111111111011, 28'b0000000000000000000000000001, 28'b1111111111111111001101100001, 28'b0000000000000000111010110111, 28'b0000000000000000001001101110, 28'b0000000000000010100101101010, 28'b1111111111111011100111010011, 28'b1111111111111111001111100111, 28'b1111111111111111110111001100, 28'b0000000000000001101110101011, 28'b1111111111111100111011010111, 28'b0000000000000000001010111000, 28'b1111111111111001111101101000, 28'b1111111111111111110110010101, 28'b1111111111111111000011000110, 28'b1111111111111111101011010111, 28'b0000000000000010010111011000, 28'b1111111111111111011001110111, 28'b1111111111111101110000000111, 28'b0000000000000000101110010000, 28'b0000000000000000000000001010, 28'b0000000000000011001010101010, 28'b0000000000000100001011111001, 28'b1111111111111101011000000010, 28'b1111111111111100011010000000}, 
{28'b0000000000000000100010100010, 28'b0000000000000000001101000100, 28'b1111111111111100101011111111, 28'b1111111111111111100010111100, 28'b1111111111111111111111111100, 28'b0000000000000000000001000111, 28'b0000000000000000110110011010, 28'b0000000000000011010010100111, 28'b0000000000000000000000000010, 28'b0000000000000000001010011000, 28'b0000000000000000100011110110, 28'b1111111111111011101011110101, 28'b1111111111111111011101111010, 28'b1111111111111011001010111000, 28'b0000000000000011110110001100, 28'b0000000000000000000000001101, 28'b1111111111111111111111100110, 28'b1111111111111010110111111010, 28'b1111111111111111111111110111, 28'b1111111111111111011001111010, 28'b1111111111111111110101010110, 28'b0000000000000000000000000000, 28'b0000000000000000011111111011, 28'b1111111111111110110011000011, 28'b0000000000000000011011001101, 28'b0000000000000011010010011000, 28'b0000000000000011011010010100, 28'b0000000000000011000111111110, 28'b0000000000000010011101101101, 28'b0000000000000000000000000110, 28'b0000000000000000111010011111, 28'b0000000000000110010001001010}, 
{28'b1111111111111111110011000101, 28'b1111111111111110000110001111, 28'b0000000000000011000111010110, 28'b1111111111111111001011010101, 28'b0000000000000000100011101110, 28'b0000000000000001010101111100, 28'b1111111111111111111111111111, 28'b1111111111111101101101000101, 28'b1111111111111111010100011000, 28'b1111111111111011001100011011, 28'b0000000000000011100101000001, 28'b0000000000000000000001111100, 28'b0000000000000011010110100100, 28'b0000000000000101010111000110, 28'b1111111111111111000100011001, 28'b1111111111111001000010001110, 28'b1111111111111111001010110101, 28'b0000000000000011110000100101, 28'b1111111111111101101111001011, 28'b1111111111111110010101001011, 28'b0000000000000000011110011011, 28'b0000000000000000000000100000, 28'b1111111111111011101000111101, 28'b1111111111111110011110000100, 28'b1111111111111111101011111001, 28'b1111111111111111000001101000, 28'b0000000000000000111001011111, 28'b0000000000000101101000001111, 28'b0000000000000001111101101101, 28'b1111111111111111111111111101, 28'b0000000000000000101001010101, 28'b0000000000000000001110001001}, 
{28'b0000000000000000010101101110, 28'b0000000000000011101000010011, 28'b0000000000000000000000000011, 28'b0000000000000010010111010011, 28'b0000000000000110101001100111, 28'b1111111111111110101000100101, 28'b1111111111111111111111111101, 28'b1111111111111111101001010101, 28'b0000000000000010010110000001, 28'b1111111111111110011101111100, 28'b1111111111111111111111010101, 28'b0000000000000010101010101010, 28'b0000000000000000000100010110, 28'b0000000000000000001110000010, 28'b1111111111110011110010001010, 28'b1111111111111111010111010110, 28'b0000000000000000000000000000, 28'b0000000000000001100110110000, 28'b1111111111111111111110010010, 28'b0000000000000010011000111001, 28'b1111111111111111111111111000, 28'b1111111111111110100111100011, 28'b1111111111111011100000010011, 28'b0000000000000001000010111111, 28'b0000000000000010010010011000, 28'b1111111111110111001000000111, 28'b1111111111111111111111111001, 28'b0000000000000000000000000101, 28'b0000000000000100010110100101, 28'b1111111111111001100101101101, 28'b0000000000000000000000111011, 28'b1111111111111111111100111000}, 
{28'b0000000000000000000100110101, 28'b1111111111111101010010000111, 28'b0000000000000000011011101000, 28'b1111111111111111111000010110, 28'b0000000000000000011010101010, 28'b0000000000000100001110111000, 28'b1111111111111010001100111011, 28'b0000000000000000010001100111, 28'b0000000000000011011000110010, 28'b1111111111111101010011010110, 28'b1111111111111111110100000111, 28'b0000000000000000011001000010, 28'b1111111111111111111011011011, 28'b0000000000000001011011100101, 28'b0000000000000000110110111110, 28'b1111111111111111110111011111, 28'b0000000000000000100010010101, 28'b0000000000000000000000001001, 28'b0000000000000000001011000011, 28'b0000000000000011000010011111, 28'b1111111111111111110001101000, 28'b1111111111111100001000000000, 28'b1111111111111011001010010011, 28'b1111111111111110011100110101, 28'b1111111111111011010001100100, 28'b0000000000000001101010100000, 28'b0000000000000100111111000110, 28'b0000000000000010111100110000, 28'b1111111111111111111010101010, 28'b1111111111111101000001001110, 28'b1111111111111101100000111001, 28'b0000000000000000011110100101}, 
{28'b0000000000000000011010100101, 28'b1111111111111100001011011101, 28'b1111111111111111110111010110, 28'b0000000000000001001101000011, 28'b1111111111111100001011000001, 28'b0000000000000001010110111001, 28'b1111111111111111111111111100, 28'b1111111111111111111111111010, 28'b1111111111111111111111111110, 28'b0000000000000000000000000111, 28'b0000000000000010000111010111, 28'b1111111111111111110111001010, 28'b0000000000000000000100111111, 28'b0000000000000000000000001000, 28'b0000000000000001000001001101, 28'b1111111111111111110111010111, 28'b0000000000000000000001011010, 28'b1111111111111111111111101001, 28'b1111111111111101011011000111, 28'b1111111111111011111101000111, 28'b1111111111111111111111101101, 28'b1111111111111011101110101010, 28'b1111111111111101100101110011, 28'b1111111111111101000001101010, 28'b0000000000000111000111111110, 28'b0000000000000000001001000000, 28'b1111111111111111101000011011, 28'b0000000000000010100010011110, 28'b0000000000000111001011100000, 28'b0000000000000011001010001011, 28'b1111111111110111100001000011, 28'b1111111111111110100001000001}, 
{28'b0000000000000011000000011100, 28'b1111111111111111111111110011, 28'b0000000000000010000000100001, 28'b1111111111111111110101110101, 28'b0000000000000011110111101011, 28'b1111111111111110110110111111, 28'b0000000000000000100100010000, 28'b0000000000000011010110001000, 28'b0000000000000010001001000110, 28'b1111111111111011110100101000, 28'b1111111111111111100000011111, 28'b0000000000000000111110111010, 28'b0000000000000000100011010011, 28'b1111111111111111111000100001, 28'b0000000000000000101011011110, 28'b0000000000000000000000001000, 28'b0000000000000010111001100010, 28'b0000000000000000010001111101, 28'b0000000000000010111111100101, 28'b1111111111111111011110011101, 28'b1111111111111110111110110011, 28'b1111111111111111011001101100, 28'b1111111111111111111111111000, 28'b0000000000000010011010100011, 28'b1111111111111110011000011001, 28'b1111111111111111111100110100, 28'b0000000000000000000000000000, 28'b0000000000000000000000001000, 28'b0000000000000000000000000100, 28'b0000000000000010010101100011, 28'b1111111111111101011011110100, 28'b1111111111111111110100000111}, 
{28'b1111111111111111111111101010, 28'b1111111111111111110000001100, 28'b1111111111111100010001111000, 28'b0000000000000010010001101010, 28'b0000000000000001110010010000, 28'b1111111111111111000111111001, 28'b1111111111111111111111111011, 28'b1111111111111110001011110100, 28'b0000000000000000000011011100, 28'b1111111111111111111111110101, 28'b1111111111111101100101101100, 28'b1111111111111110000001111000, 28'b0000000000000011110101010000, 28'b0000000000000000000000000000, 28'b1111111111111110111110100110, 28'b1111111111111111111111111110, 28'b0000000000000001101101100111, 28'b1111111111111111111111111010, 28'b1111111111111111111111111111, 28'b1111111111111110010001011011, 28'b0000000000000010100001111101, 28'b0000000000000000000000000010, 28'b0000000000000001001111111101, 28'b1111111111111111110001010101, 28'b0000000000000001010000011000, 28'b0000000000000000000001001000, 28'b0000000000000000000000000011, 28'b0000000000000001111011010001, 28'b1111111111111110011101101001, 28'b1111111111111111101000011010, 28'b0000000000000001010010001101, 28'b1111111111111111001001110011}, 
{28'b1111111111111111110111011011, 28'b1111111111111101100010000000, 28'b0000000000000100110000010101, 28'b1111111111111111011110101111, 28'b0000000000000001100100100011, 28'b1111111111111101101101100001, 28'b0000000000000000000000000010, 28'b0000000000000000010001100000, 28'b1111111111111100001010101111, 28'b1111111111111111111001011101, 28'b1111111111111111000000101000, 28'b0000000000000000011101110010, 28'b1111111111111101011000000111, 28'b0000000000000001000110100110, 28'b0000000000000001100111100100, 28'b0000000000000000111000000110, 28'b0000000000000000101011111011, 28'b1111111111111111101100100001, 28'b1111111111111010010101011010, 28'b1111111111111111111001000110, 28'b1111111111111111100010110111, 28'b0000000000000001000111100110, 28'b1111111111111111000111001000, 28'b1111111111111111111111111111, 28'b0000000000000001100101001110, 28'b1111111111111111101000101011, 28'b1111111111111111111000100110, 28'b0000000000000011000111001011, 28'b1111111111111100110100001110, 28'b1111111111111101101000111000, 28'b0000000000000010110011100111, 28'b0000000000000000010010011000}, 
{28'b0000000000000011011100101001, 28'b0000000000000001100111000100, 28'b0000000000000000000000011001, 28'b1111111111111110101110100110, 28'b1111111111111111010111110100, 28'b1111111111111111111111100100, 28'b0000000000000000000000000010, 28'b1111111111111111011100100110, 28'b1111111111111111000000011010, 28'b1111111111111111000011010101, 28'b0000000000000000000000001010, 28'b0000000000000001010001000101, 28'b0000000000000000000011010001, 28'b0000000000000000011011000100, 28'b1111111111111111101001001001, 28'b0000000000000000000010111101, 28'b1111111111111110110001011110, 28'b0000000000000000000000010011, 28'b1111111111111111110110111111, 28'b1111111111111111111111101100, 28'b0000000000000000000001001100, 28'b0000000000000000011110011011, 28'b0000000000000000110001110000, 28'b0000000000000000000000000011, 28'b0000000000000000000000001001, 28'b1111111111111011000111011011, 28'b1111111111111110011001111110, 28'b0000000000000000000011011000, 28'b0000000000000000001010011110, 28'b0000000000000000000000101011, 28'b1111111111111110100101010100, 28'b0000000000000000001010111111}, 
{28'b0000000000000001100000000100, 28'b1111111111110111101001001100, 28'b1111111111111111111111111100, 28'b1111111111111111011001011111, 28'b1111111111111110001000110001, 28'b1111111111111111111011000101, 28'b0000000000000000000000000001, 28'b0000000000000100011000011110, 28'b1111111111111111101001100100, 28'b1111111111111111110100110000, 28'b0000000000000000101010001111, 28'b1111111111111010101101101110, 28'b0000000000000000001100010010, 28'b1111111111111100011111100000, 28'b0000000000000101110001111000, 28'b1111111111111111100101001111, 28'b1111111111111110001100000011, 28'b1111111111111011100111111011, 28'b1111111111111111111010100111, 28'b1111111111111010010101100110, 28'b1111111111111001100001011100, 28'b1111111111111111111111110110, 28'b0000000000000000000000001110, 28'b0000000000000000000000000010, 28'b0000000000000001111100111100, 28'b1111111111111111111000110111, 28'b1111111111111101100111010100, 28'b1111111111111111011010110010, 28'b1111111111111111110100000100, 28'b0000000000000000000000000111, 28'b1111111111111111101111110001, 28'b1111111111111010011001101000}
};

localparam logic signed [27:0] bias [32] = '{
28'b0000000000000010000111001100,  // 0.5280959606170654
28'b0000000000000011010111011010,  // 0.8414360880851746
28'b0000000000000001100101110110,  // 0.397830605506897
28'b0000000000000001101001000111,  // 0.4105983078479767
28'b1111111111110001010111100111,  // -3.657735586166382
28'b1111111111111100011010001010,  // -0.8977976441383362
28'b0000000000000110110100100001,  // 1.7051936388015747
28'b1111111111111010111001001101,  // -1.2765135765075684
28'b1111111111111101101010100011,  // -0.5837795734405518
28'b0000000000001010110011000111,  // 2.699671983718872
28'b0000000000000000110111100100,  // 0.2170683741569519
28'b0000000000000011100001101001,  // 0.8814588785171509
28'b1111111111110101011101100111,  // -2.634300947189331
28'b1111111111111000011111011010,  // -1.877297282218933
28'b0000000000000110101001100111,  // 1.6625694036483765
28'b0000000000001010111110111101,  // 2.7459704875946045
28'b1111111111111110000101100010,  // -0.47838035225868225
28'b0000000000000110110010110100,  // 1.6984987258911133
28'b0000000000000011011010110110,  // 0.8548859357833862
28'b0000000000000100000001001010,  // 1.0045719146728516
28'b0000000000000101101011011101,  // 1.4197649955749512
28'b0000000000000011010101000111,  // 0.832463800907135
28'b0000000000000010001011000111,  // 0.5434179306030273
28'b0000000000000011101101011111,  // 0.9277304410934448
28'b1111111111111110101000010010,  // -0.3426123857498169
28'b1111111111111101110000111110,  // -0.5587119460105896
28'b1111111111111101100001000011,  // -0.6208624839782715
28'b1111111111111010111000010000,  // -1.2802538871765137
28'b0000000000000000001111001101,  // 0.05940237268805504
28'b1111111111111100101101101111,  // -0.8213341236114502
28'b0000000000000011100000110111,  // 0.8783953189849854
28'b1111111111111100001100111000   // -0.949700653553009
};
endpackage