// Width: 17
// NFRAC: 8
package dense_2_17_9;

localparam logic signed [16:0] weights [64][32] = '{ 
{17'b00000000001000100, 17'b00000000000000010, 17'b11111111111001111, 17'b11111111111111010, 17'b00000000001000010, 17'b00000000000000000, 17'b11111111111011011, 17'b11111111111111111, 17'b11111111110111001, 17'b00000000000010100, 17'b00000000000000000, 17'b11111111111111110, 17'b11111111111111111, 17'b11111111111001100, 17'b11111111111110011, 17'b11111111110111100, 17'b00000000000000000, 17'b11111111111111100, 17'b11111111111001111, 17'b11111111111010111, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111111101, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000011001, 17'b00000000001100010, 17'b00000000000101100, 17'b11111111111111111, 17'b00000000000001100, 17'b11111111110010111, 17'b00000000000000000}, 
{17'b11111111111100110, 17'b11111111111011000, 17'b11111111111011100, 17'b11111111111110001, 17'b11111111111111110, 17'b00000000000001011, 17'b11111111111000110, 17'b00000000000000001, 17'b00000000000000001, 17'b11111111111101111, 17'b00000000000100111, 17'b11111111111110100, 17'b11111111111110000, 17'b11111111111001000, 17'b00000000000000001, 17'b11111111111110011, 17'b00000000000000011, 17'b11111111111001110, 17'b00000000000101011, 17'b00000000000111010, 17'b11111111111110111, 17'b11111111111111110, 17'b11111111111111111, 17'b00000000000000110, 17'b11111111111101101, 17'b00000000001000110, 17'b00000000000111111, 17'b00000000000000010, 17'b00000000000000111, 17'b11111111110000011, 17'b00000000000000001, 17'b00000000000000000}, 
{17'b00000000000010010, 17'b11111111111100010, 17'b11111111111011110, 17'b11111111111110101, 17'b11111111111101100, 17'b11111111111101010, 17'b11111111111010000, 17'b00000000000000001, 17'b11111111111011101, 17'b00000000000000010, 17'b00000000000000000, 17'b11111111111101011, 17'b00000000000010111, 17'b11111111111101111, 17'b11111111111111111, 17'b11111111111110110, 17'b00000000000000001, 17'b00000000000011000, 17'b00000000000001111, 17'b00000000000111010, 17'b00000000000001010, 17'b11111111111101010, 17'b00000000000000000, 17'b00000000000001000, 17'b11111111111111011, 17'b00000000000110101, 17'b00000000000100110, 17'b00000000000011000, 17'b11111111111111111, 17'b11111111111011001, 17'b11111111111111100, 17'b00000000000011001}, 
{17'b00000000000100011, 17'b00000000000000100, 17'b00000000000001101, 17'b11111111111111101, 17'b11111111101111101, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000000111001, 17'b00000000000111110, 17'b11111111111111100, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000000000001, 17'b11111111111111011, 17'b00000000000110110, 17'b00000000000000000, 17'b11111111111111001, 17'b11111111111111111, 17'b11111111111010010, 17'b11111111111110000, 17'b00000000000001100, 17'b11111111111101111, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111110011, 17'b00000000000010010, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111001000, 17'b00000000001001111}, 
{17'b11111111101010001, 17'b11111111111111001, 17'b11111111111111110, 17'b00000000000000001, 17'b11111111111111001, 17'b00000000000000001, 17'b11111111111110011, 17'b11111111111011001, 17'b00000000000001101, 17'b11111111111111010, 17'b11111111111111100, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000000110101, 17'b00000000000000000, 17'b00000000001010100, 17'b11111111111111111, 17'b00000000000110111, 17'b11111111110011001, 17'b00000000000000000, 17'b11111111111100011, 17'b00000000000101011, 17'b00000000001000010, 17'b00000000000000000, 17'b00000000000001011, 17'b00000000000101001, 17'b00000000000111101, 17'b00000000000000100, 17'b11111111111111110, 17'b11111111111111111, 17'b11111111111111100, 17'b00000000000111001}, 
{17'b00000000000001110, 17'b11111111111111111, 17'b00000000000100110, 17'b11111111101011001, 17'b11111111010011111, 17'b11111111110100110, 17'b00000000001011010, 17'b11111111101100000, 17'b11111111111111111, 17'b11111111101010010, 17'b11111111101111111, 17'b11111111110101000, 17'b00000000001011010, 17'b11111111111111111, 17'b11111111111111100, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111011110, 17'b11111111111111111, 17'b11111111110000010, 17'b00000000000000000, 17'b00000000000101111, 17'b11111111111111111, 17'b00000000000000101, 17'b00000000001000100, 17'b00000000000001101, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000000110100, 17'b11111111111110111, 17'b00000000000110011}, 
{17'b11111111111110110, 17'b11111111111010111, 17'b11111111111000010, 17'b11111111111110011, 17'b11111111110110110, 17'b00000000000010000, 17'b11111111111010001, 17'b11111111111011011, 17'b11111111110010101, 17'b00000000000001100, 17'b11111111111111110, 17'b11111111111010111, 17'b00000000000011110, 17'b11111111111111101, 17'b11111111111110101, 17'b11111111101110010, 17'b11111111111111111, 17'b00000000000010101, 17'b00000000000110001, 17'b11111111111010110, 17'b11111111111011001, 17'b11111111111101111, 17'b11111111111111111, 17'b00000000000000111, 17'b11111111111110100, 17'b11111111101011010, 17'b11111111110111100, 17'b11111111111110100, 17'b00000000000000001, 17'b11111111111111010, 17'b00000000000000111, 17'b11111111111111111}, 
{17'b11111111111011000, 17'b11111111111101000, 17'b11111111111101011, 17'b11111111111000011, 17'b11111111111100010, 17'b11111111111111111, 17'b00000000000011010, 17'b11111111111101011, 17'b00000000000110011, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000000111000, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111111101101, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000000001011, 17'b11111111111010001, 17'b00000000000000011, 17'b11111111111111111, 17'b11111111111101101, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111111111}, 
{17'b11111111110000101, 17'b11111111111110001, 17'b11111111110011110, 17'b00000000000011111, 17'b00000000001111100, 17'b11111111111111111, 17'b11111111111111000, 17'b00000000000111101, 17'b11111111110001111, 17'b11111111111110100, 17'b00000000000000000, 17'b11111111111001100, 17'b11111111111111111, 17'b00000000000010011, 17'b11111111111001111, 17'b00000000011000001, 17'b11111111111111101, 17'b00000000000001011, 17'b00000000000110101, 17'b00000000000111110, 17'b00000000000000000, 17'b11111111110101010, 17'b00000000000000000, 17'b00000000001101001, 17'b11111111111010001, 17'b00000000010110010, 17'b11111111111011001, 17'b11111111111001011, 17'b11111111110000111, 17'b11111111110001001, 17'b00000000000000000, 17'b00000000000001101}, 
{17'b00000000000000000, 17'b11111111111111100, 17'b11111111111101101, 17'b00000000000000000, 17'b00000000001001110, 17'b11111111111111010, 17'b11111111111101111, 17'b00000000000010111, 17'b00000000000011001, 17'b00000000000000000, 17'b11111111111111101, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111100010, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111111110, 17'b00000000000000000, 17'b00000000000010101, 17'b00000000000000100, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000000001, 17'b00000000000001001, 17'b11111111111011110, 17'b00000000000010001, 17'b00000000000111111, 17'b11111111111111111, 17'b00000000000000001, 17'b00000000000001100, 17'b00000000000010001}, 
{17'b00000000000011000, 17'b00000000000000000, 17'b11111111111100101, 17'b11111111110111111, 17'b11111111100110100, 17'b00000000000100010, 17'b00000000000000000, 17'b11111111100101100, 17'b00000000000001001, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000000000010, 17'b00000000000000000, 17'b11111111111111011, 17'b11111111110011110, 17'b11111111111111111, 17'b00000000000111000, 17'b00000000000100000, 17'b00000000000110000, 17'b11111111110001111, 17'b11111111110100100, 17'b00000000000011110, 17'b11111111111110111, 17'b11111111111110100, 17'b00000000001011011, 17'b11111111111100111, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000000110110, 17'b11111111111111111, 17'b00000000000000001}, 
{17'b11111111111001101, 17'b11111111110000001, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000001010101, 17'b11111111110111011, 17'b11111111111000111, 17'b00000000000011101, 17'b11111111111111111, 17'b00000000000100110, 17'b00000000000010010, 17'b11111111111101100, 17'b00000000000000000, 17'b00000000000000011, 17'b11111111111111010, 17'b11111111110111111, 17'b00000000000101100, 17'b00000000000000111, 17'b00000000001001100, 17'b00000000000010110, 17'b00000000000000000, 17'b11111111111110110, 17'b00000000000100000, 17'b11111111111101001, 17'b11111111110110001, 17'b11111111111111110, 17'b00000000000101111, 17'b11111111111111111, 17'b00000000000000010, 17'b11111111111100111, 17'b00000000000100011, 17'b00000000001000110}, 
{17'b00000000000000011, 17'b00000000000000000, 17'b00000000000111000, 17'b00000000000000010, 17'b11111111111110101, 17'b00000000000101110, 17'b00000000000010111, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111011100, 17'b11111111111110010, 17'b11111111111010101, 17'b11111111111111111, 17'b00000000000001100, 17'b11111111111101110, 17'b00000000011010111, 17'b00000000000000000, 17'b11111111111100111, 17'b11111111111001111, 17'b11111111111111100, 17'b00000000000110010, 17'b00000000000100000, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000000111000, 17'b00000000001000100, 17'b00000000001111110, 17'b00000000000000010, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111111100, 17'b11111111111101101}, 
{17'b11111111111011000, 17'b00000000000001100, 17'b00000000000001010, 17'b11111111111000000, 17'b11111111110111011, 17'b00000000001111000, 17'b00000000000001100, 17'b00000000000000000, 17'b11111111111010110, 17'b11111111111101001, 17'b00000000000100001, 17'b00000000000010010, 17'b00000000000000000, 17'b11111111111101011, 17'b00000000001001001, 17'b11111111111111111, 17'b11111111111111100, 17'b00000000000000000, 17'b00000000000000011, 17'b11111111111110100, 17'b00000000000010100, 17'b00000000000000100, 17'b00000000000011101, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000010101000, 17'b11111111111110001, 17'b11111111111111010, 17'b11111111111111111, 17'b11111111111100100, 17'b11111111111110101, 17'b00000000000101101}, 
{17'b00000000000001111, 17'b00000000000010010, 17'b00000000001010011, 17'b11111111111110101, 17'b00000000000011001, 17'b00000000001011001, 17'b00000000000000000, 17'b11111111111111000, 17'b00000000000011110, 17'b11111111111100010, 17'b11111111111111111, 17'b11111111111100001, 17'b00000000000000000, 17'b00000000001100100, 17'b11111111111111011, 17'b00000000000000000, 17'b00000000000111100, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111110101111, 17'b11111111111000001, 17'b11111111111110110, 17'b11111111111111111, 17'b11111111111011010, 17'b11111111111110110, 17'b11111111111101010, 17'b11111111111001101, 17'b11111111111001001, 17'b00000000000000111, 17'b00000000000011100, 17'b11111111110011010, 17'b00000000000000000}, 
{17'b11111111110110011, 17'b00000000000000000, 17'b11111111111111100, 17'b11111111111110011, 17'b11111111111111111, 17'b00000000000100010, 17'b11111111111101100, 17'b00000000001000101, 17'b11111111110100011, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111111101000, 17'b00000000000010100, 17'b00000000000101110, 17'b11111111111111101, 17'b11111111110111111, 17'b11111111111110000, 17'b00000000000011100, 17'b00000000000010000, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000000010100, 17'b11111111111000010, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111011111}, 
{17'b11111111110101001, 17'b11111111111111110, 17'b11111111111111111, 17'b11111111111111011, 17'b11111111111111110, 17'b00000000000011011, 17'b00000000000000001, 17'b00000000000001000, 17'b00000000000001001, 17'b00000000000010000, 17'b00000000000010100, 17'b00000000000101001, 17'b00000000000000110, 17'b11111111111100111, 17'b00000000000000000, 17'b00000000001100001, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000000011100, 17'b00000000000100100, 17'b00000000000000111, 17'b00000000000001010, 17'b11111111111111000, 17'b11111111111110111, 17'b00000000000000110, 17'b11111111111101110, 17'b11111111111011111, 17'b00000000000110101, 17'b11111111111111000, 17'b00000000000001000, 17'b11111111111001111}, 
{17'b00000000000000000, 17'b11111111111111111, 17'b00000000000001001, 17'b00000000000000000, 17'b00000000011101000, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000000011100, 17'b11111111111101100, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000000100001, 17'b00000000000000000, 17'b11111111111011010, 17'b11111111111111111, 17'b11111111111101110, 17'b00000000001010011, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000010001, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000001010}, 
{17'b11111111111111111, 17'b00000000000000111, 17'b11111111111111111, 17'b00000000000001100, 17'b11111111111110100, 17'b11111111111100001, 17'b11111111111110000, 17'b00000000001000111, 17'b00000000000000000, 17'b00000000000011000, 17'b11111111111111101, 17'b00000000000010000, 17'b11111111111110111, 17'b11111111111010111, 17'b11111111111001111, 17'b00000000000000011, 17'b11111111111111111, 17'b11111111111110111, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000000010011, 17'b00000000000001001, 17'b11111111111011111, 17'b00000000000011100, 17'b11111111111010101, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111010101, 17'b00000000000000000, 17'b00000000000001011, 17'b11111111111111000}, 
{17'b11111111111111101, 17'b11111111111100110, 17'b00000000000000000, 17'b11111111111110000, 17'b00000000000110111, 17'b11111111111111111, 17'b11111111111111010, 17'b00000000000011011, 17'b11111111110011011, 17'b00000000000000000, 17'b11111111111110110, 17'b11111111111111111, 17'b00000000001011001, 17'b00000000000111010, 17'b11111111111100110, 17'b11111111111111010, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111011101, 17'b11111111111100001, 17'b00000000000100001, 17'b00000000000000000, 17'b11111111111011100, 17'b00000000000000110, 17'b11111111111101011, 17'b11111111111110111, 17'b00000000000100010, 17'b00000000000000000, 17'b11111111111000000}, 
{17'b00000000010100010, 17'b00000000001010111, 17'b11111111111000000, 17'b00000000000000000, 17'b11111111110100111, 17'b00000000000000000, 17'b00000000000111001, 17'b00000000000000111, 17'b00000000000111001, 17'b11111111111111111, 17'b11111111111011000, 17'b11111111111101011, 17'b00000000000100100, 17'b00000000000000111, 17'b11111111111100110, 17'b00000000000100001, 17'b00000000010001001, 17'b11111111111011110, 17'b11111111110110100, 17'b00000000000000000, 17'b11111111111111000, 17'b11111111111010010, 17'b11111111111111100, 17'b11111111111111111, 17'b00000000000010110, 17'b11111111110100011, 17'b00000000000010110, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000011011, 17'b11111111111111000, 17'b00000000000001111}, 
{17'b11111111111101000, 17'b11111111111001110, 17'b11111111111110110, 17'b11111111111010101, 17'b11111111111111011, 17'b00000000000001100, 17'b00000000000000000, 17'b11111111111111101, 17'b00000000000001001, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111001000, 17'b00000000000011010, 17'b00000000000010100, 17'b11111111111100101, 17'b00000000001110001, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111111110, 17'b00000000000000000, 17'b00000000001010000, 17'b11111111110000111, 17'b11111111111100100, 17'b11111111111110001, 17'b11111111111111011, 17'b00000000000110010, 17'b11111111111110010, 17'b00000000000000100, 17'b00000000001111011, 17'b11111111101111100, 17'b11111111110100010, 17'b00000000000000101}, 
{17'b00000000000000100, 17'b11111111111110000, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111101000111, 17'b11111111101100100, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111110111100, 17'b00000000000000110, 17'b00000000000000000, 17'b11111111111111000, 17'b00000000000000000, 17'b11111111111110001, 17'b11111111111110010, 17'b11111111111101110, 17'b11111111111011010, 17'b00000000001001000, 17'b00000000000000000, 17'b00000000000001011, 17'b11111111111111111, 17'b11111111111101101, 17'b00000000000000000, 17'b11111111111101001, 17'b00000000000111000, 17'b11111111101100000, 17'b00000000000111000, 17'b11111111111111111, 17'b11111111111111110, 17'b00000000000110011, 17'b11111111111111111, 17'b00000000000111100}, 
{17'b11111111111111111, 17'b00000000000000001, 17'b11111111111110100, 17'b00000000000010011, 17'b00000000000001110, 17'b11111111110101000, 17'b00000000000000000, 17'b00000000000010000, 17'b00000000010010100, 17'b11111111111111101, 17'b00000000000000000, 17'b00000000000001110, 17'b00000000001011011, 17'b11111111111110111, 17'b00000000000000011, 17'b00000000000011001, 17'b11111111111111111, 17'b00000000000000111, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111110111001, 17'b00000000000001001, 17'b00000000000010001, 17'b00000000000000101, 17'b11111111111111111, 17'b00000000000110111, 17'b00000000000000001, 17'b00000000000100000, 17'b11111111110010101, 17'b00000000000011010, 17'b00000000001100101, 17'b00000000000000001}, 
{17'b11111111110100110, 17'b00000000000110110, 17'b11111111110111101, 17'b00000000000011111, 17'b11111111111100101, 17'b00000000000000000, 17'b00000000001111111, 17'b11111111111000100, 17'b11111111110110101, 17'b00000000000101011, 17'b11111111111000110, 17'b11111111111111001, 17'b11111111111111111, 17'b00000000001011000, 17'b11111111111111111, 17'b11111111110110010, 17'b11111111111111111, 17'b00000000001110000, 17'b11111111110000111, 17'b11111111111111001, 17'b00000000001010001, 17'b11111111110100011, 17'b00000000000001101, 17'b11111111111111100, 17'b00000000001000101, 17'b11111111101111101, 17'b11111111110100011, 17'b11111111111001101, 17'b11111111111111111, 17'b00000000000011010, 17'b00000000000000110, 17'b00000000000101101}, 
{17'b11111111111101000, 17'b00000000000001101, 17'b11111111111111111, 17'b00000000000100110, 17'b11111111111110110, 17'b00000000000111010, 17'b00000000000000000, 17'b11111111111111101, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000010000101, 17'b00000000000000011, 17'b00000000000110000, 17'b00000000000000000, 17'b11111111111001001, 17'b11111111111101100, 17'b11111111111111111, 17'b11111111111111011, 17'b00000000000001010, 17'b11111111111111111, 17'b11111111111010000, 17'b11111111111111111, 17'b00000000001001011, 17'b00000000001001111, 17'b11111111111111111, 17'b11111111111111011, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111111100111}, 
{17'b11111111111101011, 17'b00000000000000000, 17'b00000000001000101, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111100010, 17'b00000000000000000, 17'b11111111100100010, 17'b00000000000110111, 17'b00000000000000011, 17'b00000000000000110, 17'b11111111110100011, 17'b00000000000000000, 17'b11111111111011100, 17'b11111111111110111, 17'b00000000000000000, 17'b00000000000000101, 17'b00000000000000000, 17'b00000000000011100, 17'b00000000000000000, 17'b11111111111111101, 17'b00000000001010100, 17'b00000000001100000, 17'b11111111111000111, 17'b11111111111011011, 17'b00000000000111111, 17'b11111111110110001, 17'b00000000000000111, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000000101111}, 
{17'b11111111111100010, 17'b11111111111111111, 17'b11111111111000010, 17'b11111111111001100, 17'b11111111111111100, 17'b11111111111011101, 17'b00000000000000000, 17'b00000000000010111, 17'b11111111111000010, 17'b11111111111101010, 17'b11111111111110011, 17'b00000000000000000, 17'b00000000000000111, 17'b11111111111111101, 17'b11111111111110000, 17'b00000000000011000, 17'b00000000000111001, 17'b00000000000100001, 17'b11111111111011110, 17'b00000000000001100, 17'b11111111111111100, 17'b11111111111111000, 17'b00000000000000101, 17'b00000000000000100, 17'b11111111111101110, 17'b00000000000010110, 17'b11111111111101000, 17'b00000000000001111, 17'b11111111111111111, 17'b11111111110110100, 17'b11111111111111001, 17'b00000000000111001}, 
{17'b11111111111111001, 17'b11111111111101010, 17'b00000000000010011, 17'b00000000001000000, 17'b00000000000010101, 17'b00000000000010101, 17'b00000000000001011, 17'b11111111111001100, 17'b11111111111001011, 17'b00000000000010001, 17'b00000000000000011, 17'b00000000000001011, 17'b00000000000000101, 17'b00000000000000001, 17'b00000000000110100, 17'b00000000000000001, 17'b11111111111110010, 17'b00000000000011010, 17'b11111111111111000, 17'b11111111111110110, 17'b00000000000011100, 17'b11111111111100000, 17'b11111111111111001, 17'b00000000000100000, 17'b00000000000000101, 17'b11111111111100100, 17'b11111111111001101, 17'b11111111111111100, 17'b11111111110111000, 17'b00000000000001111, 17'b00000000000011010, 17'b00000000000000000}, 
{17'b11111111111111100, 17'b11111111111111010, 17'b11111111111111100, 17'b11111111111110111, 17'b11111111111011110, 17'b11111111111011100, 17'b00000000000010000, 17'b00000000000000010, 17'b11111111111010001, 17'b00000000000101010, 17'b11111111111111010, 17'b11111111111111111, 17'b11111111111100011, 17'b00000000000000001, 17'b00000000000000111, 17'b11111111111110010, 17'b11111111111111011, 17'b11111111111110101, 17'b11111111111101011, 17'b00000000000000000, 17'b11111111111011100, 17'b00000000000011010, 17'b11111111111001001, 17'b00000000000000001, 17'b00000000000001010, 17'b00000000000011111, 17'b00000000000000110, 17'b00000000000000001, 17'b00000000001001010, 17'b00000000000001101, 17'b00000000000000000, 17'b00000000000010101}, 
{17'b11111111111111011, 17'b00000000001000000, 17'b11111111111111111, 17'b11111111111110111, 17'b11111111111001001, 17'b11111111111101100, 17'b00000000001101001, 17'b11111111101001111, 17'b11111111110100110, 17'b11111111111001100, 17'b11111111111000111, 17'b11111111110111111, 17'b11111111111111111, 17'b00000000001111011, 17'b11111111111111001, 17'b00000000000000000, 17'b11111111111001001, 17'b00000000001110010, 17'b11111111110010110, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111110101001, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000000001110, 17'b11111111111110001, 17'b11111111111011010, 17'b11111111111111111, 17'b00000000000101100, 17'b00000000000000000, 17'b11111111111101011, 17'b00000000000000000}, 
{17'b00000000001011110, 17'b11111111111100011, 17'b00000000000100001, 17'b11111111111110111, 17'b00000000000010011, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111101000, 17'b00000000000000000, 17'b00000000000010111, 17'b11111111111111111, 17'b11111111111110000, 17'b11111111111111111, 17'b00000000000111010, 17'b00000000000000100, 17'b00000000000001010, 17'b00000000000000110, 17'b11111111111111001, 17'b00000000000000101, 17'b00000000000000000, 17'b11111111111111101, 17'b11111111111111111, 17'b11111111110110001, 17'b11111111111111111, 17'b00000000000001110, 17'b11111111111100010, 17'b11111111111011101, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000010001110, 17'b11111111110110110, 17'b11111111111100010}, 
{17'b11111111111110100, 17'b11111111111100101, 17'b11111111111101111, 17'b00000000000001001, 17'b00000000000100011, 17'b11111111111011110, 17'b11111111111111111, 17'b11111111111000111, 17'b00000000000001111, 17'b00000000000100010, 17'b11111111111001001, 17'b11111111110111111, 17'b00000000000000110, 17'b11111111101010001, 17'b11111111111101100, 17'b11111111111100000, 17'b11111111111001101, 17'b11111111111111111, 17'b00000000000100010, 17'b00000000000000000, 17'b11111111111110100, 17'b11111111111110100, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111110000, 17'b11111111100111110, 17'b11111111101110001, 17'b11111111110111010, 17'b00000000000001110, 17'b00000000000110100, 17'b11111111111111111, 17'b00000000000111101}, 
{17'b11111111111101000, 17'b11111111111001001, 17'b00000000000101001, 17'b00000000000010011, 17'b00000000000001011, 17'b11111111111101000, 17'b11111111111110111, 17'b00000000000011001, 17'b00000000010001001, 17'b11111111111010100, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000000011110, 17'b11111111111110001, 17'b11111111111111011, 17'b11111111111111011, 17'b11111111111100110, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000111010, 17'b11111111111011101, 17'b11111111111111111, 17'b00000000000100000, 17'b11111111111111101, 17'b00000000000000000, 17'b00000000010000110, 17'b00000000001010011, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111110010100, 17'b11111111111101110, 17'b11111111111111111}, 
{17'b00000000000000011, 17'b00000000000001100, 17'b11111111111111100, 17'b00000000000000000, 17'b00000000000111011, 17'b11111111110000100, 17'b00000000000000000, 17'b11111111111100111, 17'b00000000000101111, 17'b00000000000000000, 17'b11111111111111011, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000000000001, 17'b11111111111100100, 17'b00000000001000010, 17'b11111111111111110, 17'b11111111111111100, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111111110, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000000000011, 17'b11111111110101110, 17'b00000000000001101, 17'b00000000000101110, 17'b11111111111111111, 17'b00000000000011000, 17'b11111111111111111, 17'b00000000000010011}, 
{17'b11111111111001100, 17'b00000000000000010, 17'b11111111110000100, 17'b00000000000000001, 17'b11111111111110011, 17'b11111111111110101, 17'b11111111111111111, 17'b11111111111101000, 17'b11111111111110110, 17'b11111111111101111, 17'b00000000000001100, 17'b00000000000000110, 17'b11111111111010010, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111111111101, 17'b00000000000010010, 17'b11111111111111010, 17'b11111111111111000, 17'b11111111111111000, 17'b11111111111111111, 17'b00000000001000101, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111111101, 17'b00000000001010001, 17'b00000000000110000, 17'b00000000000001000, 17'b11111111111100111, 17'b11111111111111101, 17'b00000000000010000, 17'b00000000000001110}, 
{17'b00000000000001000, 17'b00000000000001010, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111110001000, 17'b00000000000001011, 17'b00000000000000110, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111010100, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111010110, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111110100100, 17'b00000000000000010, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000100001, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000001110100, 17'b00000000001010111, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111000100, 17'b00000000000000000, 17'b11111111111111111}, 
{17'b00000000000010011, 17'b00000000000001101, 17'b00000000001000000, 17'b11111111111000000, 17'b00000000000100001, 17'b00000000000011110, 17'b00000000000000001, 17'b00000000000110001, 17'b00000000000000011, 17'b11111111111111100, 17'b00000000000001001, 17'b00000000000000001, 17'b11111111111111111, 17'b00000000000011110, 17'b11111111111111110, 17'b11111111111110101, 17'b00000000000000000, 17'b00000000000001000, 17'b11111111111110011, 17'b00000000000011001, 17'b00000000000001000, 17'b11111111101101011, 17'b11111111111100010, 17'b00000000000010111, 17'b11111111111111111, 17'b11111111101111110, 17'b11111111111011111, 17'b11111111111111010, 17'b11111111111111111, 17'b11111111111110001, 17'b00000000000000000, 17'b11111111111110101}, 
{17'b00000000000000000, 17'b11111111111111111, 17'b11111111111101000, 17'b11111111111010100, 17'b00000000000001010, 17'b00000000000000000, 17'b00000000000011000, 17'b11111111111111110, 17'b00000000000111111, 17'b11111111111111110, 17'b00000000000000000, 17'b11111111110101000, 17'b11111111111111111, 17'b00000000000100000, 17'b11111111111111111, 17'b11111111110111101, 17'b00000000000000000, 17'b11111111111111101, 17'b00000000001000011, 17'b11111111111111111, 17'b11111111110010000, 17'b11111111111111111, 17'b00000000001000010, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000000100011, 17'b11111111111100111, 17'b00000000000010001, 17'b00000000000000000, 17'b11111111111001100, 17'b00000000000000000, 17'b00000000000000000}, 
{17'b11111111111001000, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111111110, 17'b00000000001111110, 17'b11111111111100000, 17'b11111111111111110, 17'b11111111111111110, 17'b11111111111110100, 17'b11111111111110011, 17'b00000000000010000, 17'b00000000000100010, 17'b11111111111110110, 17'b00000000000111111, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111110110111, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111101011, 17'b00000000000000000, 17'b00000000000001001, 17'b00000000000000011, 17'b11111111111111101, 17'b11111111111110010, 17'b11111111111001100, 17'b11111111110110100, 17'b00000000000000000, 17'b11111111111100011, 17'b00000000000001010, 17'b11111111111111111, 17'b00000000000010011}, 
{17'b11111111110010110, 17'b11111111111010111, 17'b11111111111011000, 17'b00000000000000000, 17'b00000000010010010, 17'b11111111111000111, 17'b00000000000000000, 17'b11111111111110010, 17'b11111111110010111, 17'b00000000000100011, 17'b11111111111111111, 17'b00000000010010001, 17'b00000000000000000, 17'b11111111111110011, 17'b11111111111111111, 17'b00000000000001000, 17'b11111111111111011, 17'b00000000000000000, 17'b11111111111110100, 17'b00000000001111110, 17'b00000000000001001, 17'b11111111111110101, 17'b00000000000011100, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111100111, 17'b11111111111110100, 17'b11111111110001000, 17'b11111111111011011, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111110000}, 
{17'b00000000000111001, 17'b11111111100110011, 17'b11111111101000110, 17'b11111111111010100, 17'b00000000010101011, 17'b11111111111111111, 17'b11111111110100111, 17'b00000000001000011, 17'b00000000000001111, 17'b00000000000000000, 17'b00000000000110101, 17'b11111111110111010, 17'b00000000000000000, 17'b00000000000000001, 17'b11111111111110111, 17'b00000000000000100, 17'b11111111111100101, 17'b11111111100010100, 17'b00000000000101010, 17'b00000000001011000, 17'b00000000001000011, 17'b00000000000000000, 17'b00000000000000111, 17'b11111111110011000, 17'b11111111101011110, 17'b11111111111111110, 17'b11111111110110011, 17'b11111111110001010, 17'b11111111111001110, 17'b11111111100011111, 17'b00000000001101011, 17'b00000000001101101}, 
{17'b00000000000000000, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000001000010, 17'b11111111111010000, 17'b00000000000000100, 17'b00000000000010010, 17'b11111111110100110, 17'b00000000000001001, 17'b11111111111111110, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000000111101, 17'b00000000000001101, 17'b00000000000000101, 17'b00000000000001111, 17'b00000000001010101, 17'b11111111111001000, 17'b00000000000000000, 17'b11111111111010101, 17'b11111111111111111, 17'b00000000001010000, 17'b00000000000000010, 17'b11111111111111111, 17'b11111111101110000, 17'b11111111111111101, 17'b11111111111011000, 17'b11111111111110000, 17'b00000000000000000, 17'b00000000000100010, 17'b00000000000011010}, 
{17'b11111111111110100, 17'b00000000000100010, 17'b11111111110110010, 17'b00000000000000101, 17'b00000000000110001, 17'b11111111111110101, 17'b11111111111111110, 17'b00000000000101001, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111111101111, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111110111, 17'b11111111111100000, 17'b11111111111101111, 17'b11111111111110001, 17'b11111111111101111, 17'b11111111111100011, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111111110100, 17'b11111111111101110, 17'b00000000001100101, 17'b00000000000000000, 17'b11111111110100011, 17'b11111111111111101, 17'b00000000000011111, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000001000000, 17'b11111111111111111}, 
{17'b11111111111111111, 17'b00000000000000001, 17'b11111111111111111, 17'b11111111111011000, 17'b11111111100100011, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111111110, 17'b11111111101100110, 17'b00000000000010100, 17'b11111111111100110, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111110100001, 17'b11111111111110100, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000000010, 17'b00000000000001001, 17'b00000000001011000, 17'b11111111111100001, 17'b11111111110110011, 17'b00000000000000000, 17'b11111111110111101, 17'b11111111111100110, 17'b11111111111000100, 17'b11111111111111110, 17'b11111111111111100, 17'b11111111111111011, 17'b11111111110000111, 17'b11111111111110111, 17'b00000000000111110}, 
{17'b00000000000011100, 17'b00000000000111000, 17'b11111111111111111, 17'b00000000000101000, 17'b11111111111001010, 17'b11111111111100000, 17'b00000000000011000, 17'b00000000000010001, 17'b11111111111110011, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111110101101, 17'b11111111111111111, 17'b00000000000100100, 17'b11111111111100010, 17'b00000000000001000, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000000110101, 17'b11111111110101100, 17'b00000000001000111, 17'b00000000000001100, 17'b00000000000000000, 17'b00000000000110110, 17'b00000000000000000, 17'b11111111111110110, 17'b11111111110011110, 17'b11111111111100011, 17'b11111111111010100, 17'b00000000000101101}, 
{17'b00000000000000000, 17'b00000000000000001, 17'b11111111110100010, 17'b11111111111111111, 17'b00000000000110100, 17'b11111111111011011, 17'b11111111111111100, 17'b11111111111111111, 17'b00000000000000101, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111001011, 17'b00000000000011000, 17'b00000000000000001, 17'b00000000000000000, 17'b00000000000001001, 17'b11111111111111111, 17'b11111111111011001, 17'b00000000000000100, 17'b00000000000000000, 17'b11111111111110111, 17'b11111111111111010, 17'b00000000001001011, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111110110101, 17'b11111111110101100, 17'b00000000000111101, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000000000111, 17'b00000000001001000}, 
{17'b11111111110101000, 17'b11111111111111111, 17'b11111111111001001, 17'b00000000000000001, 17'b11111111110100101, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111111101111, 17'b11111111101110111, 17'b11111111111111001, 17'b00000000000000000, 17'b11111111111111101, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111111101, 17'b11111111111110011, 17'b11111111111011010, 17'b11111111111100111, 17'b00000000000010000, 17'b11111111111111111, 17'b11111111111111001, 17'b00000000000000000, 17'b00000000001010110, 17'b11111111111111111, 17'b00000000000100110, 17'b00000000000010111, 17'b11111111111011100, 17'b00000000000110110, 17'b11111111111110100, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000010010101}, 
{17'b11111111110101111, 17'b00000000000000111, 17'b00000000000001100, 17'b11111111111111000, 17'b00000000000111110, 17'b11111111110110010, 17'b11111111111111110, 17'b00000000001000011, 17'b00000000000101000, 17'b00000000000000010, 17'b11111111111111111, 17'b11111111111101110, 17'b11111111111101001, 17'b11111111111101111, 17'b11111111111110011, 17'b00000000000010111, 17'b11111111111111111, 17'b00000000000000010, 17'b00000000000100100, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000000000011, 17'b00000000001000000, 17'b00000000000001011, 17'b00000000000000001, 17'b11111111111100100, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111111100, 17'b11111111111111100, 17'b11111111111111111, 17'b00000000000010001}, 
{17'b11111111111111111, 17'b00000000000000000, 17'b11111111111001001, 17'b11111111111101100, 17'b00000000001001000, 17'b11111111111111111, 17'b11111111111101100, 17'b00000000000111110, 17'b11111111111110010, 17'b00000000001001010, 17'b00000000000010101, 17'b11111111111100001, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111111100, 17'b00000000000000101, 17'b11111111111101100, 17'b11111111110111100, 17'b00000000001000111, 17'b00000000000100111, 17'b00000000010100010, 17'b00000000000110011, 17'b00000000000111111, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000000001110, 17'b00000000000010100, 17'b11111111110010100, 17'b11111111111111111, 17'b11111111111111110, 17'b11111111111111110}, 
{17'b00000000000000000, 17'b11111111111101001, 17'b11111111111100101, 17'b00000000000000000, 17'b11111111111000001, 17'b00000000000000000, 17'b00000000000110001, 17'b00000000000011011, 17'b00000000000001101, 17'b11111111111100110, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111110101, 17'b00000000000110011, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111110110010, 17'b00000000000000000, 17'b11111111111001110, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111111110, 17'b00000000000000011, 17'b00000000000000100, 17'b00000000000000111, 17'b00000000000100011, 17'b11111111111101111, 17'b11111111111111110, 17'b11111111110001101, 17'b00000000000010100}, 
{17'b00000000001110001, 17'b11111111111111101, 17'b00000000000010000, 17'b11111111111100101, 17'b11111111111101010, 17'b00000000000001000, 17'b00000000000101001, 17'b00000000000000000, 17'b00000000010000110, 17'b00000000000000000, 17'b11111111111111010, 17'b00000000000000100, 17'b00000000000011000, 17'b11111111111111111, 17'b00000000000001101, 17'b00000000000011010, 17'b11111111111111110, 17'b11111111110001110, 17'b11111111111110001, 17'b11111111111111111, 17'b00000000000011101, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000000011100, 17'b00000000000000100, 17'b11111111110111100, 17'b11111111111100101, 17'b00000000000100001, 17'b11111111111111000, 17'b00000000001000010, 17'b11111111111111111, 17'b11111111111010010}, 
{17'b00000000000000011, 17'b00000000000011010, 17'b11111111111111111, 17'b11111111111110110, 17'b11111111110100101, 17'b11111111111111111, 17'b00000000000001011, 17'b11111111111110100, 17'b00000000000101010, 17'b11111111111110111, 17'b11111111111111111, 17'b11111111111110111, 17'b11111111111111111, 17'b11111111111110110, 17'b00000000000000000, 17'b00000000001010000, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000000001000, 17'b00000000000100000, 17'b00000000000000000, 17'b00000000000000001, 17'b00000000000001000, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000000101, 17'b00000000000000000, 17'b00000000000011000}, 
{17'b11111111110110000, 17'b00000000000100001, 17'b00000000000000100, 17'b11111111111100101, 17'b11111111110011001, 17'b11111111111111011, 17'b00000000000010001, 17'b11111111110011010, 17'b00000000010000010, 17'b00000000000010010, 17'b00000000000000100, 17'b00000000000011000, 17'b00000000000001011, 17'b00000000000000000, 17'b00000000001101000, 17'b11111111111101010, 17'b00000000000000001, 17'b00000000000000000, 17'b11111111111111110, 17'b00000000000000000, 17'b11111111110010001, 17'b00000000000000100, 17'b00000000000100111, 17'b00000000000001001, 17'b00000000000001001, 17'b11111111101010111, 17'b11111111110101000, 17'b11111111111000010, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000001010011, 17'b11111111111001011}, 
{17'b11111111111111100, 17'b11111111111001110, 17'b11111111111100101, 17'b11111111110010111, 17'b11111111110111101, 17'b00000000001010110, 17'b00000000001001111, 17'b11111111111010100, 17'b00000000000001010, 17'b11111111111110110, 17'b11111111111100111, 17'b11111111110111111, 17'b00000000000011010, 17'b11111111110110111, 17'b00000000000110000, 17'b11111111111111111, 17'b00000000001010101, 17'b11111111111111111, 17'b11111111111111110, 17'b11111111111011101, 17'b11111111111110101, 17'b11111111111101111, 17'b11111111110111011, 17'b00000000000010101, 17'b11111111111111111, 17'b11111111111111110, 17'b11111111111000101, 17'b00000000001010000, 17'b00000000001000111, 17'b11111111111101000, 17'b11111111101011110, 17'b00000000000100100}, 
{17'b00000000000000000, 17'b11111111111111001, 17'b11111111111111111, 17'b11111111111100111, 17'b00000000000000111, 17'b00000000000000010, 17'b00000000000010001, 17'b00000000000000001, 17'b00000000000011110, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000011000, 17'b00000000000000000, 17'b00000000000000011, 17'b11111111111011110, 17'b11111111111100100, 17'b00000000000000000, 17'b00000000000101110, 17'b00000000000001110, 17'b00000000000100000, 17'b11111111111111011, 17'b11111111111010111, 17'b11111111111111111, 17'b00000000000010011, 17'b11111111111111111, 17'b00000000000001000, 17'b11111111111111110, 17'b00000000000010001, 17'b00000000000000000, 17'b00000000000010101, 17'b11111111110011110, 17'b11111111111111111}, 
{17'b00000000001001111, 17'b11111111111111101, 17'b00000000000100110, 17'b11111111110110001, 17'b11111111111001110, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000000000111, 17'b00000000000000000, 17'b11111111111011111, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111011110, 17'b00000000000100100, 17'b11111111111111111, 17'b11111111111111000, 17'b00000000000000000, 17'b00000000000011110, 17'b11111111111001100, 17'b00000000000011101, 17'b00000000000100011, 17'b00000000000100001, 17'b11111111111111111, 17'b00000000010001101, 17'b11111111111011000, 17'b00000000001011101, 17'b11111111111110010, 17'b11111111110100011, 17'b11111111111010011, 17'b00000000000100011}, 
{17'b11111111101110100, 17'b11111111111111001, 17'b11111111111011000, 17'b11111111111111111, 17'b00000000001000010, 17'b11111111111010010, 17'b11111111111110000, 17'b00000000000111100, 17'b00000000000011000, 17'b11111111111000011, 17'b00000000000000000, 17'b11111111111111000, 17'b11111111111111101, 17'b00000000000100011, 17'b11111111111000001, 17'b11111111111111101, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111111111011, 17'b00000000000000000, 17'b11111111111001111, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111110101011, 17'b00000000000010001, 17'b00000000010011110, 17'b00000000001011000, 17'b11111111111110110, 17'b11111111111010110, 17'b11111111110001101, 17'b00000000000000000, 17'b11111111111110011}, 
{17'b00000000000000101, 17'b00000000000110110, 17'b00000000000000101, 17'b11111111111011001, 17'b00000000000000001, 17'b11111111111111001, 17'b00000000000000000, 17'b00000000000110101, 17'b00000000000110111, 17'b11111111111011101, 17'b00000000000100011, 17'b00000000000000110, 17'b11111111111111111, 17'b11111111111111100, 17'b11111111111010111, 17'b00000000001000000, 17'b11111111111110101, 17'b11111111110101101, 17'b00000000000011101, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000000011101, 17'b11111111111101100, 17'b11111111111111110, 17'b11111111111110010, 17'b00000000000010110, 17'b11111111111011100, 17'b00000000000100010, 17'b11111111110100010, 17'b00000000000010100, 17'b11111111111111111, 17'b00000000000101000}, 
{17'b11111111111110101, 17'b00000000000000000, 17'b00000000000010110, 17'b00000000000000000, 17'b11111111111110000, 17'b11111111111111111, 17'b00000000000011010, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000000001, 17'b00000000000000000, 17'b00000000000000101, 17'b11111111111100100, 17'b00000000000000010, 17'b00000000000011100, 17'b00000000000001011, 17'b00000000000011011, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000000100000, 17'b00000000000111111, 17'b11111111111100110, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000000000010, 17'b11111111110001001, 17'b11111111111111111, 17'b11111111111101101, 17'b11111111111111111, 17'b00000000010010000, 17'b00000000000000000, 17'b11111111111001011}, 
{17'b11111111111111001, 17'b11111111111100001, 17'b11111111111111101, 17'b00000000000000001, 17'b00000000000010111, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111111010, 17'b00000000000010010, 17'b11111111111111101, 17'b00000000000000000, 17'b00000000000001000, 17'b00000000001001011, 17'b11111111111100101, 17'b00000000000000011, 17'b11111111100100110, 17'b11111111111111101, 17'b11111111111110000, 17'b00000000000000010, 17'b11111111111110011, 17'b00000000000010111, 17'b11111111111000110, 17'b00000000000011101, 17'b00000000000011010, 17'b11111111111111100, 17'b11111111101001001, 17'b11111111111000101, 17'b11111111111111010, 17'b11111111111111011, 17'b00000000001100011, 17'b11111111111111110, 17'b00000000000100111}, 
{17'b00000000000001100, 17'b00000000000000000, 17'b00000000000101100, 17'b11111111111100010, 17'b11111111111101110, 17'b00000000000111100, 17'b11111111111010111, 17'b00000000000001110, 17'b11111111110110000, 17'b00000000000000010, 17'b00000000000000100, 17'b11111111111101010, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111001111, 17'b00000000001101110, 17'b11111111111000000, 17'b11111111111111100, 17'b00000000000011110, 17'b11111111111111111, 17'b00000000000010001, 17'b11111111110000101, 17'b00000000001010000, 17'b11111111111111111, 17'b11111111111100000, 17'b00000000001111100, 17'b00000000000100101, 17'b11111111111010111, 17'b11111111111011101, 17'b11111111101110110, 17'b11111111111111101, 17'b00000000000000100}, 
{17'b11111111111111111, 17'b00000000000000001, 17'b11111111111110111, 17'b11111111110111011, 17'b11111111111111111, 17'b11111111110011011, 17'b00000000000000000, 17'b00000000001001101, 17'b00000000000111110, 17'b00000000000000100, 17'b00000000000000000, 17'b11111111111100011, 17'b00000000001010101, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000001101111, 17'b00000000000000000, 17'b11111111111110101, 17'b11111111111110010, 17'b11111111110101101, 17'b00000000000100001, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000000001000, 17'b11111111111101101, 17'b11111111110001010, 17'b00000000001000110, 17'b11111111110001110, 17'b00000000000001101, 17'b11111111111101011, 17'b00000000000000000}, 
{17'b00000000000001111, 17'b00000000000101111, 17'b00000000000000010, 17'b11111111111111111, 17'b11111111110001010, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000000111110, 17'b00000000001000110, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000000101011, 17'b11111111111100101, 17'b11111111110010001, 17'b11111111111110111, 17'b11111111111100110, 17'b11111111111100111, 17'b11111111111101110, 17'b11111111111111111, 17'b11111111111101111, 17'b11111111111111010, 17'b11111111111111101, 17'b00000000000100100, 17'b11111111111111111, 17'b00000000001110110}
};

localparam logic signed [16:0] bias [32] = '{
17'b00000000101111001,  // 1.474280834197998
17'b00000000010110001,  // 0.6914801001548767
17'b00000000101110000,  // 1.4406442642211914
17'b00000000101101000,  // 1.408045768737793
17'b00000000011111100,  // 0.9864811301231384
17'b00000000011011101,  // 0.8636202812194824
17'b11111111101100010,  // -0.6153604388237
17'b00000000001111011,  // 0.4839226007461548
17'b00000000001111100,  // 0.4862793982028961
17'b00000000001011111,  // 0.37162142992019653
17'b00000000001110101,  // 0.45989668369293213
17'b00000000101001100,  // 1.2998151779174805
17'b11111111011111011,  // -1.016528844833374
17'b11111111110100101,  // -0.35249894857406616
17'b00000000001110010,  // 0.44582197070121765
17'b11111111111100011,  // -0.1119980737566948
17'b11111111111101110,  // -0.06717441976070404
17'b00000000000000001,  // 0.00487547367811203
17'b00000000000110001,  // 0.1946917623281479
17'b11111111100111000,  // -0.7796769738197327
17'b00000000010111010,  // 0.7287401556968689
17'b00000000110110111,  // 1.714877724647522
17'b11111111001100111,  // -1.5971007347106934
17'b00000000000010010,  // 0.07393483817577362
17'b00000000001010010,  // 0.3225609362125397
17'b00000000011011000,  // 0.8453295230865479
17'b00000000011100110,  // 0.898597240447998
17'b00000000001000001,  // 0.2548799514770508
17'b00000000011111001,  // 0.9735668301582336
17'b00000000100100000,  // 1.1261906623840332
17'b00000000001110010,  // 0.44768181443214417
17'b11111110110100001   // -2.3676068782806396
};
endpackage