// Width: 18
// NFRAC: 9
package dense_4_18_9;

localparam logic signed [17:0] weights [32][5] = '{ 
{18'b111111111111111001, 18'b000000000010100001, 18'b111111111101100111, 18'b000000000000100001, 18'b111111111111001001}, 
{18'b111111111011100010, 18'b111111111111100011, 18'b000000000011101011, 18'b111111111111111001, 18'b000000000000001000}, 
{18'b000000000010111110, 18'b000000000001101100, 18'b111111111111110001, 18'b111111111100110000, 18'b111111111110010100}, 
{18'b111111111100111111, 18'b111111111101000001, 18'b111111111111000110, 18'b000000000010011101, 18'b000000000001111000}, 
{18'b000000000000111110, 18'b000000000001000001, 18'b000000000001010000, 18'b111111111111110110, 18'b111111110111111001}, 
{18'b000000000010100111, 18'b111111111100110110, 18'b000000000001011100, 18'b111111111110101101, 18'b111111111110101000}, 
{18'b111111111100110010, 18'b000000000000010010, 18'b111111111111111111, 18'b000000000001011001, 18'b000000000000100011}, 
{18'b111111111111111111, 18'b000000000010010001, 18'b111111111100110111, 18'b000000000001010011, 18'b000000000001000101}, 
{18'b000000000001010011, 18'b111111111110101001, 18'b000000000000000000, 18'b111111111100010011, 18'b111111111110000000}, 
{18'b111111111111111111, 18'b111111111101110111, 18'b000000000001011011, 18'b000000000011011100, 18'b000000000000000000}, 
{18'b111111111110111101, 18'b111111111110110101, 18'b000000000000000000, 18'b000000000100101001, 18'b111111111101110110}, 
{18'b000000000001010110, 18'b000000000001110101, 18'b111111111101010001, 18'b111111111111110001, 18'b000000000000111110}, 
{18'b000000000000000000, 18'b000000000001010101, 18'b000000000000000100, 18'b111111111110010101, 18'b111111111011000001}, 
{18'b000000000001011010, 18'b000000000000100000, 18'b000000000011010110, 18'b111111111111011100, 18'b111111111100100100}, 
{18'b000000000000101110, 18'b111111111111100111, 18'b111111111101000111, 18'b111111111111101111, 18'b000000000100010010}, 
{18'b111111111100001101, 18'b111111111110000010, 18'b111111111110001110, 18'b000000000011001100, 18'b000000000000010000}, 
{18'b000000000010110001, 18'b111111111110101000, 18'b111111111110111010, 18'b111111111110001100, 18'b111111111111100001}, 
{18'b000000000001100011, 18'b111111111111101011, 18'b111111111100101100, 18'b111111111111110000, 18'b000000000000100100}, 
{18'b000000000010000100, 18'b000000000000010101, 18'b111111111110010000, 18'b000000000000000000, 18'b111111111100111111}, 
{18'b000000000001110110, 18'b111111111111010011, 18'b111111111110010011, 18'b000000000001101010, 18'b000000000000110000}, 
{18'b000000000000100010, 18'b111111111111110000, 18'b000000000010011000, 18'b111111111100100011, 18'b111111111111110101}, 
{18'b000000000000000000, 18'b000000000000111100, 18'b000000000011111001, 18'b111111111011110110, 18'b111111111011000011}, 
{18'b111111111111001101, 18'b000000000000111000, 18'b000000000001011010, 18'b111111111101001001, 18'b000000000100001011}, 
{18'b111111111111111111, 18'b000000000001010100, 18'b000000000010010000, 18'b000000000000010011, 18'b111111111011011011}, 
{18'b111111111110101001, 18'b000000000010111010, 18'b111111111110001101, 18'b000000000000000010, 18'b000000000011000110}, 
{18'b000000000000001101, 18'b000000000010001000, 18'b000000000000001111, 18'b111111111010000001, 18'b000000000100011000}, 
{18'b111111111100010100, 18'b111111111110000011, 18'b000000000001101101, 18'b000000000001111101, 18'b000000000001100111}, 
{18'b000000000000000010, 18'b000000000001111011, 18'b111111111111101101, 18'b111111111110110010, 18'b000000000000010000}, 
{18'b111111111111001010, 18'b000000000001111110, 18'b111111111011111110, 18'b000000000001000111, 18'b111111111110101110}, 
{18'b111111111111110110, 18'b000000000001001000, 18'b111111111110101001, 18'b111111111100110010, 18'b000000000100101111}, 
{18'b000000000011100101, 18'b000000000000100011, 18'b000000000010100110, 18'b111111111011010010, 18'b111111111101011110}, 
{18'b111111111111100001, 18'b111111111100111010, 18'b000000000010111011, 18'b000000000000100100, 18'b000000000001000001}
};

localparam logic signed [17:0] bias [5] = '{
18'b111111111111100000,  // -0.06223141402006149
18'b111111111111011111,  // -0.06270556896924973
18'b111111111111011100,  // -0.07014333456754684
18'b000000000000101010,  // 0.0820775106549263
18'b000000000001101110   // 0.2155742198228836
};
endpackage