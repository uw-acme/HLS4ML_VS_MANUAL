// Width: 8
// NFRAC: 4
package dense_2_8_4;

localparam logic signed [7:0] weights [64][32] = '{ 
{8'b00000100, 8'b00000000, 8'b11111100, 8'b11111111, 8'b00000100, 8'b00000000, 8'b11111101, 8'b11111111, 8'b11111011, 8'b00000001, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111100, 8'b11111111, 8'b11111011, 8'b00000000, 8'b11111111, 8'b11111100, 8'b11111101, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000001, 8'b00000110, 8'b00000010, 8'b11111111, 8'b00000000, 8'b11111001, 8'b00000000}, 
{8'b11111110, 8'b11111101, 8'b11111101, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111100, 8'b00000000, 8'b00000000, 8'b11111110, 8'b00000010, 8'b11111111, 8'b11111111, 8'b11111100, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111100, 8'b00000010, 8'b00000011, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111110, 8'b00000100, 8'b00000011, 8'b00000000, 8'b00000000, 8'b11111000, 8'b00000000, 8'b00000000}, 
{8'b00000001, 8'b11111110, 8'b11111101, 8'b11111111, 8'b11111110, 8'b11111110, 8'b11111101, 8'b00000000, 8'b11111101, 8'b00000000, 8'b00000000, 8'b11111110, 8'b00000001, 8'b11111110, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000001, 8'b00000000, 8'b00000011, 8'b00000000, 8'b11111110, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000011, 8'b00000010, 8'b00000001, 8'b11111111, 8'b11111101, 8'b11111111, 8'b00000001}, 
{8'b00000010, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11110111, 8'b00000000, 8'b00000000, 8'b00000011, 8'b00000011, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000011, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111101, 8'b11111111, 8'b00000000, 8'b11111110, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000001, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111100, 8'b00000100}, 
{8'b11110101, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111111, 8'b11111101, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000011, 8'b00000000, 8'b00000101, 8'b11111111, 8'b00000011, 8'b11111001, 8'b00000000, 8'b11111110, 8'b00000010, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000011}, 
{8'b00000000, 8'b11111111, 8'b00000010, 8'b11110101, 8'b11101001, 8'b11111010, 8'b00000101, 8'b11110110, 8'b11111111, 8'b11110101, 8'b11110111, 8'b11111010, 8'b00000101, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111101, 8'b11111111, 8'b11111000, 8'b00000000, 8'b00000010, 8'b11111111, 8'b00000000, 8'b00000100, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000011, 8'b11111111, 8'b00000011}, 
{8'b11111111, 8'b11111101, 8'b11111100, 8'b11111111, 8'b11111011, 8'b00000001, 8'b11111101, 8'b11111101, 8'b11111001, 8'b00000000, 8'b11111111, 8'b11111101, 8'b00000001, 8'b11111111, 8'b11111111, 8'b11110111, 8'b11111111, 8'b00000001, 8'b00000011, 8'b11111101, 8'b11111101, 8'b11111110, 8'b11111111, 8'b00000000, 8'b11111111, 8'b11110101, 8'b11111011, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111111}, 
{8'b11111101, 8'b11111110, 8'b11111110, 8'b11111100, 8'b11111110, 8'b11111111, 8'b00000001, 8'b11111110, 8'b00000011, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000011, 8'b00000000, 8'b11111111, 8'b11111110, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111101, 8'b00000000, 8'b11111111, 8'b11111110, 8'b11111111, 8'b00000000, 8'b11111111}, 
{8'b11111000, 8'b11111111, 8'b11111001, 8'b00000001, 8'b00000111, 8'b11111111, 8'b11111111, 8'b00000011, 8'b11111000, 8'b11111111, 8'b00000000, 8'b11111100, 8'b11111111, 8'b00000001, 8'b11111100, 8'b00001100, 8'b11111111, 8'b00000000, 8'b00000011, 8'b00000011, 8'b00000000, 8'b11111010, 8'b00000000, 8'b00000110, 8'b11111101, 8'b00001011, 8'b11111101, 8'b11111100, 8'b11111000, 8'b11111000, 8'b00000000, 8'b00000000}, 
{8'b00000000, 8'b11111111, 8'b11111110, 8'b00000000, 8'b00000100, 8'b11111111, 8'b11111110, 8'b00000001, 8'b00000001, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111110, 8'b11111111, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000001, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111101, 8'b00000001, 8'b00000011, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000001}, 
{8'b00000001, 8'b00000000, 8'b11111110, 8'b11111011, 8'b11110011, 8'b00000010, 8'b00000000, 8'b11110010, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111001, 8'b11111111, 8'b00000011, 8'b00000010, 8'b00000011, 8'b11111000, 8'b11111010, 8'b00000001, 8'b11111111, 8'b11111111, 8'b00000101, 8'b11111110, 8'b11111111, 8'b11111111, 8'b00000011, 8'b11111111, 8'b00000000}, 
{8'b11111100, 8'b11111000, 8'b00000000, 8'b11111111, 8'b00000101, 8'b11111011, 8'b11111100, 8'b00000001, 8'b11111111, 8'b00000010, 8'b00000001, 8'b11111110, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111011, 8'b00000010, 8'b00000000, 8'b00000100, 8'b00000001, 8'b00000000, 8'b11111111, 8'b00000010, 8'b11111110, 8'b11111011, 8'b11111111, 8'b00000010, 8'b11111111, 8'b00000000, 8'b11111110, 8'b00000010, 8'b00000100}, 
{8'b00000000, 8'b00000000, 8'b00000011, 8'b00000000, 8'b11111111, 8'b00000010, 8'b00000001, 8'b11111111, 8'b00000000, 8'b11111101, 8'b11111111, 8'b11111101, 8'b11111111, 8'b00000000, 8'b11111110, 8'b00001101, 8'b00000000, 8'b11111110, 8'b11111100, 8'b11111111, 8'b00000011, 8'b00000010, 8'b00000000, 8'b11111111, 8'b00000011, 8'b00000100, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111110}, 
{8'b11111101, 8'b00000000, 8'b00000000, 8'b11111100, 8'b11111011, 8'b00000111, 8'b00000000, 8'b00000000, 8'b11111101, 8'b11111110, 8'b00000010, 8'b00000001, 8'b00000000, 8'b11111110, 8'b00000100, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000001, 8'b00000000, 8'b00000001, 8'b11111111, 8'b00000000, 8'b00001010, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111110, 8'b11111111, 8'b00000010}, 
{8'b00000000, 8'b00000001, 8'b00000101, 8'b11111111, 8'b00000001, 8'b00000101, 8'b00000000, 8'b11111111, 8'b00000001, 8'b11111110, 8'b11111111, 8'b11111110, 8'b00000000, 8'b00000110, 8'b11111111, 8'b00000000, 8'b00000011, 8'b00000000, 8'b00000000, 8'b11111010, 8'b11111100, 8'b11111111, 8'b11111111, 8'b11111101, 8'b11111111, 8'b11111110, 8'b11111100, 8'b11111100, 8'b00000000, 8'b00000001, 8'b11111001, 8'b00000000}, 
{8'b11111011, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000010, 8'b11111110, 8'b00000100, 8'b11111010, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111110, 8'b00000001, 8'b00000010, 8'b11111111, 8'b11111011, 8'b11111111, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000001, 8'b11111100, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000000, 8'b11111101}, 
{8'b11111010, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000010, 8'b00000000, 8'b11111110, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000001, 8'b00000010, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111110, 8'b11111101, 8'b00000011, 8'b11111111, 8'b00000000, 8'b11111100}, 
{8'b00000000, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00001110, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000001, 8'b11111110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000000, 8'b11111101, 8'b11111111, 8'b11111110, 8'b00000101, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000001, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000}, 
{8'b11111111, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111111, 8'b11111110, 8'b11111111, 8'b00000100, 8'b00000000, 8'b00000001, 8'b11111111, 8'b00000001, 8'b11111111, 8'b11111101, 8'b11111100, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000001, 8'b00000000, 8'b11111101, 8'b00000001, 8'b11111101, 8'b00000000, 8'b00000000, 8'b11111101, 8'b00000000, 8'b00000000, 8'b11111111}, 
{8'b11111111, 8'b11111110, 8'b00000000, 8'b11111111, 8'b00000011, 8'b11111111, 8'b11111111, 8'b00000001, 8'b11111001, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000101, 8'b00000011, 8'b11111110, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000000, 8'b11111101, 8'b11111110, 8'b00000010, 8'b00000000, 8'b11111101, 8'b00000000, 8'b11111110, 8'b11111111, 8'b00000010, 8'b00000000, 8'b11111100}, 
{8'b00001010, 8'b00000101, 8'b11111100, 8'b00000000, 8'b11111010, 8'b00000000, 8'b00000011, 8'b00000000, 8'b00000011, 8'b11111111, 8'b11111101, 8'b11111110, 8'b00000010, 8'b00000000, 8'b11111110, 8'b00000010, 8'b00001000, 8'b11111101, 8'b11111011, 8'b00000000, 8'b11111111, 8'b11111101, 8'b11111111, 8'b11111111, 8'b00000001, 8'b11111010, 8'b00000001, 8'b11111111, 8'b00000000, 8'b00000001, 8'b11111111, 8'b00000000}, 
{8'b11111110, 8'b11111100, 8'b11111111, 8'b11111101, 8'b11111111, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111100, 8'b00000001, 8'b00000001, 8'b11111110, 8'b00000111, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000101, 8'b11111000, 8'b11111110, 8'b11111111, 8'b11111111, 8'b00000011, 8'b11111111, 8'b00000000, 8'b00000111, 8'b11110111, 8'b11111010, 8'b00000000}, 
{8'b00000000, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11110100, 8'b11110110, 8'b00000000, 8'b11111111, 8'b11111011, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111110, 8'b11111101, 8'b00000100, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111110, 8'b00000000, 8'b11111110, 8'b00000011, 8'b11110110, 8'b00000011, 8'b11111111, 8'b11111111, 8'b00000011, 8'b11111111, 8'b00000011}, 
{8'b11111111, 8'b00000000, 8'b11111111, 8'b00000001, 8'b00000000, 8'b11111010, 8'b00000000, 8'b00000001, 8'b00001001, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000101, 8'b11111111, 8'b00000000, 8'b00000001, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111011, 8'b00000000, 8'b00000001, 8'b00000000, 8'b11111111, 8'b00000011, 8'b00000000, 8'b00000010, 8'b11111001, 8'b00000001, 8'b00000110, 8'b00000000}, 
{8'b11111010, 8'b00000011, 8'b11111011, 8'b00000001, 8'b11111110, 8'b00000000, 8'b00000111, 8'b11111100, 8'b11111011, 8'b00000010, 8'b11111100, 8'b11111111, 8'b11111111, 8'b00000101, 8'b11111111, 8'b11111011, 8'b11111111, 8'b00000111, 8'b11111000, 8'b11111111, 8'b00000101, 8'b11111010, 8'b00000000, 8'b11111111, 8'b00000100, 8'b11110111, 8'b11111010, 8'b11111100, 8'b11111111, 8'b00000001, 8'b00000000, 8'b00000010}, 
{8'b11111110, 8'b00000000, 8'b11111111, 8'b00000010, 8'b11111111, 8'b00000011, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00001000, 8'b00000000, 8'b00000011, 8'b00000000, 8'b11111100, 8'b11111110, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111111, 8'b11111101, 8'b11111111, 8'b00000100, 8'b00000100, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111111, 8'b11111110}, 
{8'b11111110, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000000, 8'b11111110, 8'b00000000, 8'b11110010, 8'b00000011, 8'b00000000, 8'b00000000, 8'b11111010, 8'b00000000, 8'b11111101, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000000, 8'b11111111, 8'b00000101, 8'b00000110, 8'b11111100, 8'b11111101, 8'b00000011, 8'b11111011, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000010}, 
{8'b11111110, 8'b11111111, 8'b11111100, 8'b11111100, 8'b11111111, 8'b11111101, 8'b00000000, 8'b00000001, 8'b11111100, 8'b11111110, 8'b11111111, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000001, 8'b00000011, 8'b00000010, 8'b11111101, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b11111110, 8'b00000001, 8'b11111110, 8'b00000000, 8'b11111111, 8'b11111011, 8'b11111111, 8'b00000011}, 
{8'b11111111, 8'b11111110, 8'b00000001, 8'b00000100, 8'b00000001, 8'b00000001, 8'b00000000, 8'b11111100, 8'b11111100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b00000000, 8'b11111111, 8'b00000001, 8'b11111111, 8'b11111111, 8'b00000001, 8'b11111110, 8'b11111111, 8'b00000010, 8'b00000000, 8'b11111110, 8'b11111100, 8'b11111111, 8'b11111011, 8'b00000000, 8'b00000001, 8'b00000000}, 
{8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111101, 8'b11111101, 8'b00000001, 8'b00000000, 8'b11111101, 8'b00000010, 8'b11111111, 8'b11111111, 8'b11111110, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111110, 8'b00000000, 8'b11111101, 8'b00000001, 8'b11111100, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000001}, 
{8'b11111111, 8'b00000100, 8'b11111111, 8'b11111111, 8'b11111100, 8'b11111110, 8'b00000110, 8'b11110100, 8'b11111010, 8'b11111100, 8'b11111100, 8'b11111011, 8'b11111111, 8'b00000111, 8'b11111111, 8'b00000000, 8'b11111100, 8'b00000111, 8'b11111001, 8'b00000000, 8'b11111111, 8'b11111010, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111111, 8'b11111101, 8'b11111111, 8'b00000010, 8'b00000000, 8'b11111110, 8'b00000000}, 
{8'b00000101, 8'b11111110, 8'b00000010, 8'b11111111, 8'b00000001, 8'b11111111, 8'b11111111, 8'b11111110, 8'b00000000, 8'b00000001, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000011, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111011, 8'b11111111, 8'b00000000, 8'b11111110, 8'b11111101, 8'b11111111, 8'b11111111, 8'b00001000, 8'b11111011, 8'b11111110}, 
{8'b11111111, 8'b11111110, 8'b11111110, 8'b00000000, 8'b00000010, 8'b11111101, 8'b11111111, 8'b11111100, 8'b00000000, 8'b00000010, 8'b11111100, 8'b11111011, 8'b00000000, 8'b11110101, 8'b11111110, 8'b11111110, 8'b11111100, 8'b11111111, 8'b00000010, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11110011, 8'b11110111, 8'b11111011, 8'b00000000, 8'b00000011, 8'b11111111, 8'b00000011}, 
{8'b11111110, 8'b11111100, 8'b00000010, 8'b00000001, 8'b00000000, 8'b11111110, 8'b11111111, 8'b00000001, 8'b00001000, 8'b11111101, 8'b11111111, 8'b11111111, 8'b00000001, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111110, 8'b11111111, 8'b00000000, 8'b00000011, 8'b11111101, 8'b11111111, 8'b00000010, 8'b11111111, 8'b00000000, 8'b00001000, 8'b00000101, 8'b00000000, 8'b00000000, 8'b11111001, 8'b11111110, 8'b11111111}, 
{8'b00000000, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000011, 8'b11111000, 8'b00000000, 8'b11111110, 8'b00000010, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111110, 8'b00000100, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111010, 8'b00000000, 8'b00000010, 8'b11111111, 8'b00000001, 8'b11111111, 8'b00000001}, 
{8'b11111100, 8'b00000000, 8'b11111000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111110, 8'b11111111, 8'b11111110, 8'b00000000, 8'b00000000, 8'b11111101, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000001, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000100, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000101, 8'b00000011, 8'b00000000, 8'b11111110, 8'b11111111, 8'b00000001, 8'b00000000}, 
{8'b00000000, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111101, 8'b11111111, 8'b00000000, 8'b11111101, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111010, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000010, 8'b11111111, 8'b00000000, 8'b00000111, 8'b00000101, 8'b00000000, 8'b00000000, 8'b11111100, 8'b00000000, 8'b11111111}, 
{8'b00000001, 8'b00000000, 8'b00000100, 8'b11111100, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000011, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000001, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000001, 8'b00000000, 8'b11110110, 8'b11111110, 8'b00000001, 8'b11111111, 8'b11110111, 8'b11111101, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111111}, 
{8'b00000000, 8'b11111111, 8'b11111110, 8'b11111101, 8'b00000000, 8'b00000000, 8'b00000001, 8'b11111111, 8'b00000011, 8'b11111111, 8'b00000000, 8'b11111010, 8'b11111111, 8'b00000010, 8'b11111111, 8'b11111011, 8'b00000000, 8'b11111111, 8'b00000100, 8'b11111111, 8'b11111001, 8'b11111111, 8'b00000100, 8'b11111111, 8'b11111111, 8'b00000010, 8'b11111110, 8'b00000001, 8'b00000000, 8'b11111100, 8'b00000000, 8'b00000000}, 
{8'b11111100, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000111, 8'b11111110, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000001, 8'b00000010, 8'b11111111, 8'b00000011, 8'b00000000, 8'b11111111, 8'b11111011, 8'b11111111, 8'b00000000, 8'b11111110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111100, 8'b11111011, 8'b00000000, 8'b11111110, 8'b00000000, 8'b11111111, 8'b00000001}, 
{8'b11111001, 8'b11111101, 8'b11111101, 8'b00000000, 8'b00001001, 8'b11111100, 8'b00000000, 8'b11111111, 8'b11111001, 8'b00000010, 8'b11111111, 8'b00001001, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000111, 8'b00000000, 8'b11111111, 8'b00000001, 8'b11111111, 8'b11111111, 8'b11111110, 8'b11111111, 8'b11111000, 8'b11111101, 8'b11111111, 8'b11111111, 8'b11111111}, 
{8'b00000011, 8'b11110011, 8'b11110100, 8'b11111101, 8'b00001010, 8'b11111111, 8'b11111010, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11111011, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111110, 8'b11110001, 8'b00000010, 8'b00000101, 8'b00000100, 8'b00000000, 8'b00000000, 8'b11111001, 8'b11110101, 8'b11111111, 8'b11111011, 8'b11111000, 8'b11111100, 8'b11110001, 8'b00000110, 8'b00000110}, 
{8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000100, 8'b11111101, 8'b00000000, 8'b00000001, 8'b11111010, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000011, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000101, 8'b11111100, 8'b00000000, 8'b11111101, 8'b11111111, 8'b00000101, 8'b00000000, 8'b11111111, 8'b11110111, 8'b11111111, 8'b11111101, 8'b11111111, 8'b00000000, 8'b00000010, 8'b00000001}, 
{8'b11111111, 8'b00000010, 8'b11111011, 8'b00000000, 8'b00000011, 8'b11111111, 8'b11111111, 8'b00000010, 8'b00000000, 8'b11111111, 8'b11111110, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111110, 8'b11111110, 8'b11111111, 8'b11111110, 8'b11111110, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111110, 8'b00000110, 8'b00000000, 8'b11111010, 8'b11111111, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000100, 8'b11111111}, 
{8'b11111111, 8'b00000000, 8'b11111111, 8'b11111101, 8'b11110010, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11110110, 8'b00000001, 8'b11111110, 8'b11111111, 8'b00000000, 8'b11111010, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000101, 8'b11111110, 8'b11111011, 8'b00000000, 8'b11111011, 8'b11111110, 8'b11111100, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111000, 8'b11111111, 8'b00000011}, 
{8'b00000001, 8'b00000011, 8'b11111111, 8'b00000010, 8'b11111100, 8'b11111110, 8'b00000001, 8'b00000001, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111010, 8'b11111111, 8'b00000010, 8'b11111110, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000011, 8'b11111010, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b00000000, 8'b11111111, 8'b11111001, 8'b11111110, 8'b11111101, 8'b00000010}, 
{8'b00000000, 8'b00000000, 8'b11111010, 8'b11111111, 8'b00000011, 8'b11111101, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111101, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000100, 8'b11111111, 8'b00000000, 8'b11111011, 8'b11111010, 8'b00000011, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000100}, 
{8'b11111010, 8'b11111111, 8'b11111100, 8'b00000000, 8'b11111010, 8'b00000000, 8'b11111111, 8'b11111110, 8'b11110111, 8'b11111111, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111101, 8'b11111110, 8'b00000001, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000101, 8'b11111111, 8'b00000010, 8'b00000001, 8'b11111101, 8'b00000011, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00001001}, 
{8'b11111010, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000011, 8'b11111011, 8'b11111111, 8'b00000100, 8'b00000010, 8'b00000000, 8'b11111111, 8'b11111110, 8'b11111110, 8'b11111110, 8'b11111111, 8'b00000001, 8'b11111111, 8'b00000000, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000000, 8'b11111110, 8'b11111111, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000001}, 
{8'b11111111, 8'b00000000, 8'b11111100, 8'b11111110, 8'b00000100, 8'b11111111, 8'b11111110, 8'b00000011, 8'b11111111, 8'b00000100, 8'b00000001, 8'b11111110, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111110, 8'b11111011, 8'b00000100, 8'b00000010, 8'b00001010, 8'b00000011, 8'b00000011, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b11111001, 8'b11111111, 8'b11111111, 8'b11111111}, 
{8'b00000000, 8'b11111110, 8'b11111110, 8'b00000000, 8'b11111100, 8'b00000000, 8'b00000011, 8'b00000001, 8'b00000000, 8'b11111110, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000011, 8'b11111111, 8'b11111111, 8'b11111011, 8'b00000000, 8'b11111100, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b11111110, 8'b11111111, 8'b11111000, 8'b00000001}, 
{8'b00000111, 8'b11111111, 8'b00000001, 8'b11111110, 8'b11111110, 8'b00000000, 8'b00000010, 8'b00000000, 8'b00001000, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000001, 8'b11111111, 8'b00000000, 8'b00000001, 8'b11111111, 8'b11111000, 8'b11111111, 8'b11111111, 8'b00000001, 8'b00000000, 8'b11111111, 8'b00000001, 8'b00000000, 8'b11111011, 8'b11111110, 8'b00000010, 8'b11111111, 8'b00000100, 8'b11111111, 8'b11111101}, 
{8'b00000000, 8'b00000001, 8'b11111111, 8'b11111111, 8'b11111010, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000010, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000101, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001}, 
{8'b11111011, 8'b00000010, 8'b00000000, 8'b11111110, 8'b11111001, 8'b11111111, 8'b00000001, 8'b11111001, 8'b00001000, 8'b00000001, 8'b00000000, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000110, 8'b11111110, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111001, 8'b00000000, 8'b00000010, 8'b00000000, 8'b00000000, 8'b11110101, 8'b11111010, 8'b11111100, 8'b00000000, 8'b11111111, 8'b00000101, 8'b11111100}, 
{8'b11111111, 8'b11111100, 8'b11111110, 8'b11111001, 8'b11111011, 8'b00000101, 8'b00000100, 8'b11111101, 8'b00000000, 8'b11111111, 8'b11111110, 8'b11111011, 8'b00000001, 8'b11111011, 8'b00000011, 8'b11111111, 8'b00000101, 8'b11111111, 8'b11111111, 8'b11111101, 8'b11111111, 8'b11111110, 8'b11111011, 8'b00000001, 8'b11111111, 8'b11111111, 8'b11111100, 8'b00000101, 8'b00000100, 8'b11111110, 8'b11110101, 8'b00000010}, 
{8'b00000000, 8'b11111111, 8'b11111111, 8'b11111110, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000000, 8'b00000001, 8'b11111111, 8'b00000000, 8'b00000001, 8'b00000000, 8'b00000000, 8'b11111101, 8'b11111110, 8'b00000000, 8'b00000010, 8'b00000000, 8'b00000010, 8'b11111111, 8'b11111101, 8'b11111111, 8'b00000001, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000001, 8'b00000000, 8'b00000001, 8'b11111001, 8'b11111111}, 
{8'b00000100, 8'b11111111, 8'b00000010, 8'b11111011, 8'b11111100, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b11111101, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111101, 8'b00000010, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000001, 8'b11111100, 8'b00000001, 8'b00000010, 8'b00000010, 8'b11111111, 8'b00001000, 8'b11111101, 8'b00000101, 8'b11111111, 8'b11111010, 8'b11111101, 8'b00000010}, 
{8'b11110111, 8'b11111111, 8'b11111101, 8'b11111111, 8'b00000100, 8'b11111101, 8'b11111111, 8'b00000011, 8'b00000001, 8'b11111100, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000010, 8'b11111100, 8'b11111111, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111100, 8'b11111111, 8'b00000000, 8'b11111010, 8'b00000001, 8'b00001001, 8'b00000101, 8'b11111111, 8'b11111101, 8'b11111000, 8'b00000000, 8'b11111111}, 
{8'b00000000, 8'b00000011, 8'b00000000, 8'b11111101, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000011, 8'b00000011, 8'b11111101, 8'b00000010, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111101, 8'b00000100, 8'b11111111, 8'b11111010, 8'b00000001, 8'b11111111, 8'b11111111, 8'b00000001, 8'b11111110, 8'b11111111, 8'b11111111, 8'b00000001, 8'b11111101, 8'b00000010, 8'b11111010, 8'b00000001, 8'b11111111, 8'b00000010}, 
{8'b11111111, 8'b00000000, 8'b00000001, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000001, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111110, 8'b00000000, 8'b00000001, 8'b00000000, 8'b00000001, 8'b11111111, 8'b11111111, 8'b00000010, 8'b00000011, 8'b11111110, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111000, 8'b11111111, 8'b11111110, 8'b11111111, 8'b00001001, 8'b00000000, 8'b11111100}, 
{8'b11111111, 8'b11111110, 8'b11111111, 8'b00000000, 8'b00000001, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000001, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000100, 8'b11111110, 8'b00000000, 8'b11110010, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000001, 8'b11111100, 8'b00000001, 8'b00000001, 8'b11111111, 8'b11110100, 8'b11111100, 8'b11111111, 8'b11111111, 8'b00000110, 8'b11111111, 8'b00000010}, 
{8'b00000000, 8'b00000000, 8'b00000010, 8'b11111110, 8'b11111110, 8'b00000011, 8'b11111101, 8'b00000000, 8'b11111011, 8'b00000000, 8'b00000000, 8'b11111110, 8'b00000000, 8'b00000000, 8'b11111100, 8'b00000110, 8'b11111100, 8'b11111111, 8'b00000001, 8'b11111111, 8'b00000001, 8'b11111000, 8'b00000101, 8'b11111111, 8'b11111110, 8'b00000111, 8'b00000010, 8'b11111101, 8'b11111101, 8'b11110111, 8'b11111111, 8'b00000000}, 
{8'b11111111, 8'b00000000, 8'b11111111, 8'b11111011, 8'b11111111, 8'b11111001, 8'b00000000, 8'b00000100, 8'b00000011, 8'b00000000, 8'b00000000, 8'b11111110, 8'b00000101, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000110, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111010, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111110, 8'b11111000, 8'b00000100, 8'b11111000, 8'b00000000, 8'b11111110, 8'b00000000}, 
{8'b00000000, 8'b00000010, 8'b00000000, 8'b11111111, 8'b11111000, 8'b00000000, 8'b11111111, 8'b00000011, 8'b00000100, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000010, 8'b11111110, 8'b11111001, 8'b11111111, 8'b11111110, 8'b11111110, 8'b11111110, 8'b11111111, 8'b11111110, 8'b11111111, 8'b11111111, 8'b00000010, 8'b11111111, 8'b00000111}
};

localparam logic signed [7:0] bias [32] = '{
8'b00010111,  // 1.474280834197998
8'b00001011,  // 0.6914801001548767
8'b00010111,  // 1.4406442642211914
8'b00010110,  // 1.408045768737793
8'b00001111,  // 0.9864811301231384
8'b00001101,  // 0.8636202812194824
8'b11110110,  // -0.6153604388237
8'b00000111,  // 0.4839226007461548
8'b00000111,  // 0.4862793982028961
8'b00000101,  // 0.37162142992019653
8'b00000111,  // 0.45989668369293213
8'b00010100,  // 1.2998151779174805
8'b11101111,  // -1.016528844833374
8'b11111010,  // -0.35249894857406616
8'b00000111,  // 0.44582197070121765
8'b11111110,  // -0.1119980737566948
8'b11111110,  // -0.06717441976070404
8'b00000000,  // 0.00487547367811203
8'b00000011,  // 0.1946917623281479
8'b11110011,  // -0.7796769738197327
8'b00001011,  // 0.7287401556968689
8'b00011011,  // 1.714877724647522
8'b11100110,  // -1.5971007347106934
8'b00000001,  // 0.07393483817577362
8'b00000101,  // 0.3225609362125397
8'b00001101,  // 0.8453295230865479
8'b00001110,  // 0.898597240447998
8'b00000100,  // 0.2548799514770508
8'b00001111,  // 0.9735668301582336
8'b00010010,  // 1.1261906623840332
8'b00000111,  // 0.44768181443214417
8'b11011010   // -2.3676068782806396
};
endpackage