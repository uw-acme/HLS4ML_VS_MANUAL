// Width: 20
// NFRAC: 10
package dense_4_20_10;

localparam logic signed [19:0] weights [32][5] = '{ 
{20'b11111111111111110011, 20'b00000000000101000011, 20'b11111111111011001110, 20'b00000000000001000011, 20'b11111111111110010011}, 
{20'b11111111110111000100, 20'b11111111111111000111, 20'b00000000000111010111, 20'b11111111111111110011, 20'b00000000000000010001}, 
{20'b00000000000101111100, 20'b00000000000011011000, 20'b11111111111111100011, 20'b11111111111001100000, 20'b11111111111100101000}, 
{20'b11111111111001111111, 20'b11111111111010000010, 20'b11111111111110001101, 20'b00000000000100111011, 20'b00000000000011110000}, 
{20'b00000000000001111101, 20'b00000000000010000011, 20'b00000000000010100000, 20'b11111111111111101101, 20'b11111111101111110010}, 
{20'b00000000000101001110, 20'b11111111111001101100, 20'b00000000000010111001, 20'b11111111111101011010, 20'b11111111111101010001}, 
{20'b11111111111001100101, 20'b00000000000000100100, 20'b11111111111111111111, 20'b00000000000010110010, 20'b00000000000001000110}, 
{20'b11111111111111111110, 20'b00000000000100100011, 20'b11111111111001101110, 20'b00000000000010100110, 20'b00000000000010001011}, 
{20'b00000000000010100111, 20'b11111111111101010010, 20'b00000000000000000001, 20'b11111111111000100111, 20'b11111111111100000001}, 
{20'b11111111111111111111, 20'b11111111111011101111, 20'b00000000000010110110, 20'b00000000000110111000, 20'b00000000000000000000}, 
{20'b11111111111101111010, 20'b11111111111101101011, 20'b00000000000000000000, 20'b00000000001001010011, 20'b11111111111011101101}, 
{20'b00000000000010101101, 20'b00000000000011101010, 20'b11111111111010100011, 20'b11111111111111100011, 20'b00000000000001111100}, 
{20'b00000000000000000000, 20'b00000000000010101011, 20'b00000000000000001001, 20'b11111111111100101011, 20'b11111111110110000010}, 
{20'b00000000000010110101, 20'b00000000000001000001, 20'b00000000000110101101, 20'b11111111111110111000, 20'b11111111111001001001}, 
{20'b00000000000001011100, 20'b11111111111111001110, 20'b11111111111010001110, 20'b11111111111111011110, 20'b00000000001000100101}, 
{20'b11111111111000011010, 20'b11111111111100000101, 20'b11111111111100011100, 20'b00000000000110011000, 20'b00000000000000100000}, 
{20'b00000000000101100010, 20'b11111111111101010000, 20'b11111111111101110101, 20'b11111111111100011000, 20'b11111111111111000010}, 
{20'b00000000000011000111, 20'b11111111111111010110, 20'b11111111111001011001, 20'b11111111111111100000, 20'b00000000000001001000}, 
{20'b00000000000100001000, 20'b00000000000000101010, 20'b11111111111100100000, 20'b00000000000000000000, 20'b11111111111001111111}, 
{20'b00000000000011101100, 20'b11111111111110100111, 20'b11111111111100100110, 20'b00000000000011010100, 20'b00000000000001100001}, 
{20'b00000000000001000101, 20'b11111111111111100000, 20'b00000000000100110000, 20'b11111111111001000110, 20'b11111111111111101010}, 
{20'b00000000000000000000, 20'b00000000000001111000, 20'b00000000000111110010, 20'b11111111110111101101, 20'b11111111110110000111}, 
{20'b11111111111110011011, 20'b00000000000001110000, 20'b00000000000010110101, 20'b11111111111010010010, 20'b00000000001000010110}, 
{20'b11111111111111111111, 20'b00000000000010101000, 20'b00000000000100100001, 20'b00000000000000100110, 20'b11111111110110110110}, 
{20'b11111111111101010010, 20'b00000000000101110101, 20'b11111111111100011011, 20'b00000000000000000101, 20'b00000000000110001101}, 
{20'b00000000000000011010, 20'b00000000000100010000, 20'b00000000000000011110, 20'b11111111110100000010, 20'b00000000001000110001}, 
{20'b11111111111000101001, 20'b11111111111100000110, 20'b00000000000011011011, 20'b00000000000011111010, 20'b00000000000011001110}, 
{20'b00000000000000000100, 20'b00000000000011110110, 20'b11111111111111011010, 20'b11111111111101100101, 20'b00000000000000100000}, 
{20'b11111111111110010101, 20'b00000000000011111100, 20'b11111111110111111100, 20'b00000000000010001110, 20'b11111111111101011101}, 
{20'b11111111111111101101, 20'b00000000000010010000, 20'b11111111111101010011, 20'b11111111111001100101, 20'b00000000001001011111}, 
{20'b00000000000111001011, 20'b00000000000001000111, 20'b00000000000101001100, 20'b11111111110110100100, 20'b11111111111010111101}, 
{20'b11111111111111000011, 20'b11111111111001110100, 20'b00000000000101110110, 20'b00000000000001001000, 20'b00000000000010000010}
};

localparam logic signed [19:0] bias [5] = '{
20'b11111111111111000000,  // -0.06223141402006149
20'b11111111111110111111,  // -0.06270556896924973
20'b11111111111110111000,  // -0.07014333456754684
20'b00000000000001010100,  // 0.0820775106549263
20'b00000000000011011100   // 0.2155742198228836
};
endpackage