// Width: 9
// NFRAC: 4
package dense_1_9_4;

localparam logic signed [8:0] weights [16][64] = '{ 
{9'b000000100, 9'b111110101, 9'b111111101, 9'b111111100, 9'b111111001, 9'b000000001, 9'b111101111, 9'b000000000, 9'b000000000, 9'b000000100, 9'b000000000, 9'b111111001, 9'b111111111, 9'b000000011, 9'b000000000, 9'b111111011, 9'b000000011, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000110, 9'b111111010, 9'b111111111, 9'b000000111, 9'b111111010, 9'b111110101, 9'b111111011, 9'b111111100, 9'b111111110, 9'b111111111, 9'b000000000, 9'b000000011, 9'b000000011, 9'b111111111, 9'b000000000, 9'b000000100, 9'b111111111, 9'b111111011, 9'b000000000, 9'b000000011, 9'b111111111, 9'b000000100, 9'b111111011, 9'b000001110, 9'b111111111, 9'b000000111, 9'b000000000, 9'b000000010, 9'b000000011, 9'b111111111, 9'b000000000, 9'b000000010, 9'b000000011, 9'b000000001, 9'b111111110, 9'b111111011, 9'b000001000, 9'b111111000, 9'b000000111, 9'b111111010, 9'b000001100, 9'b111111111, 9'b000000000, 9'b000000001}, 
{9'b000000000, 9'b111111010, 9'b111111101, 9'b111111011, 9'b111111010, 9'b000000001, 9'b111110011, 9'b111111111, 9'b111111100, 9'b000000010, 9'b000000000, 9'b111111110, 9'b000000011, 9'b000000000, 9'b111111111, 9'b000000011, 9'b111111111, 9'b000000000, 9'b111111101, 9'b111111011, 9'b000000111, 9'b111111110, 9'b000000000, 9'b000001011, 9'b000000100, 9'b111111100, 9'b111111100, 9'b111111111, 9'b111111110, 9'b111111001, 9'b111111111, 9'b000000111, 9'b000000100, 9'b000001000, 9'b000001010, 9'b000000000, 9'b111111110, 9'b111111001, 9'b000000000, 9'b000000011, 9'b000000000, 9'b000000011, 9'b111111100, 9'b000000100, 9'b000000010, 9'b000000000, 9'b111111010, 9'b000000001, 9'b000000100, 9'b000000000, 9'b000000000, 9'b000010010, 9'b111111110, 9'b111111110, 9'b111111111, 9'b111111111, 9'b000000100, 9'b111111010, 9'b000001111, 9'b000000000, 9'b000001000, 9'b000000011, 9'b000001101, 9'b000000010}, 
{9'b111111111, 9'b000000000, 9'b111111110, 9'b111111101, 9'b111111101, 9'b000000000, 9'b000010111, 9'b111111111, 9'b111101011, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111100, 9'b000000000, 9'b111111111, 9'b000000010, 9'b000001110, 9'b111111111, 9'b000000001, 9'b000000000, 9'b000000110, 9'b111110100, 9'b000001001, 9'b111110100, 9'b000001111, 9'b111111010, 9'b111111100, 9'b111110100, 9'b000010100, 9'b000000100, 9'b000000000, 9'b000001000, 9'b000010000, 9'b111101100, 9'b111111110, 9'b000000000, 9'b111111100, 9'b000001110, 9'b111111111, 9'b000000101, 9'b000000101, 9'b000000101, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000010, 9'b111111011, 9'b111111101, 9'b111111111, 9'b000000110, 9'b111111101, 9'b000000010, 9'b111111111, 9'b000000010, 9'b111111101, 9'b111111111, 9'b111111011, 9'b111110101, 9'b111111111, 9'b000000000, 9'b000011000, 9'b000000000, 9'b111111111, 9'b111111011}, 
{9'b111111000, 9'b111111010, 9'b111110100, 9'b000000100, 9'b111111010, 9'b111101010, 9'b111111110, 9'b111111011, 9'b000000011, 9'b111111111, 9'b000010100, 9'b111111110, 9'b111110011, 9'b000001001, 9'b000000000, 9'b111111111, 9'b111111000, 9'b111111111, 9'b000000000, 9'b111111100, 9'b111101101, 9'b111111110, 9'b111110100, 9'b000000011, 9'b111111001, 9'b111110001, 9'b000000101, 9'b000001011, 9'b000010100, 9'b111111000, 9'b111110110, 9'b000000001, 9'b000001000, 9'b111110010, 9'b111111010, 9'b000000000, 9'b111110100, 9'b000000011, 9'b111111000, 9'b000000001, 9'b000000111, 9'b000000010, 9'b000000000, 9'b000000000, 9'b000001000, 9'b111111100, 9'b111111111, 9'b111111010, 9'b111111111, 9'b111111110, 9'b111110110, 9'b000000001, 9'b111111111, 9'b000000011, 9'b000000101, 9'b000001010, 9'b111110000, 9'b111110001, 9'b111110100, 9'b000001101, 9'b000011011, 9'b111110001, 9'b111111111, 9'b000000110}, 
{9'b000000101, 9'b111110110, 9'b111111011, 9'b111111111, 9'b111111101, 9'b000000101, 9'b000000011, 9'b111111111, 9'b111110110, 9'b111111100, 9'b111111010, 9'b000000000, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000101, 9'b000000010, 9'b111111001, 9'b000000000, 9'b000000000, 9'b000000011, 9'b111111110, 9'b000000001, 9'b111111111, 9'b000010001, 9'b111111101, 9'b111111011, 9'b111111001, 9'b000000000, 9'b000000010, 9'b000000001, 9'b000000100, 9'b111111111, 9'b000000001, 9'b000000010, 9'b111111111, 9'b000000000, 9'b000001110, 9'b111111011, 9'b111111110, 9'b000000110, 9'b000000011, 9'b111111000, 9'b000000000, 9'b111101110, 9'b111111111, 9'b111111110, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000011, 9'b111111111, 9'b000000101, 9'b111111100, 9'b111110100, 9'b111111000, 9'b111110111, 9'b111110110, 9'b000001011, 9'b000010101, 9'b000001100, 9'b000000001, 9'b111111111}, 
{9'b111111000, 9'b111110101, 9'b000000000, 9'b000000100, 9'b000000100, 9'b111111100, 9'b000001001, 9'b111111111, 9'b000000011, 9'b111111111, 9'b111111111, 9'b111111110, 9'b111111101, 9'b000001001, 9'b111111110, 9'b000000000, 9'b111110110, 9'b111111010, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111010, 9'b111111010, 9'b000000111, 9'b111111010, 9'b111111111, 9'b000000100, 9'b111111110, 9'b111110001, 9'b111111111, 9'b111111110, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000010, 9'b000000101, 9'b000000000, 9'b111111110, 9'b111111011, 9'b111111111, 9'b111111101, 9'b111110111, 9'b000000110, 9'b000000000, 9'b000001001, 9'b000000000, 9'b111111111, 9'b000000001, 9'b111111001, 9'b000000011, 9'b000000000, 9'b111111110, 9'b111111010, 9'b000000110, 9'b111111111, 9'b000000101, 9'b000000011, 9'b000000011, 9'b111111111, 9'b111111111, 9'b111110011, 9'b111111101, 9'b111111111, 9'b111111111}, 
{9'b111111011, 9'b111111010, 9'b111111001, 9'b111111110, 9'b111111101, 9'b000000001, 9'b111110100, 9'b111111101, 9'b111111100, 9'b111111111, 9'b111111011, 9'b000000101, 9'b000000000, 9'b000000010, 9'b000000100, 9'b000000000, 9'b000001100, 9'b000000001, 9'b000000011, 9'b000000100, 9'b111111101, 9'b000000101, 9'b111111100, 9'b111110111, 9'b000000010, 9'b000001000, 9'b111111111, 9'b000000000, 9'b111110000, 9'b000000100, 9'b000000100, 9'b111111010, 9'b000000111, 9'b000001010, 9'b000000000, 9'b000000101, 9'b111111111, 9'b000000100, 9'b000000011, 9'b000000000, 9'b111111110, 9'b111111010, 9'b000000010, 9'b000000111, 9'b000001000, 9'b111111101, 9'b111111110, 9'b111111100, 9'b111111101, 9'b000000001, 9'b000000000, 9'b000000000, 9'b000000000, 9'b000000010, 9'b111111101, 9'b000001100, 9'b000000101, 9'b111111111, 9'b000000110, 9'b000000011, 9'b111100101, 9'b111110110, 9'b111111101, 9'b111111111}, 
{9'b000000000, 9'b000000011, 9'b111111111, 9'b111111111, 9'b111111010, 9'b111111111, 9'b111111011, 9'b000000000, 9'b000000000, 9'b000000110, 9'b000000000, 9'b111111001, 9'b111111110, 9'b000000000, 9'b111111111, 9'b111111000, 9'b111110010, 9'b111111111, 9'b111110110, 9'b111111000, 9'b111111001, 9'b000000101, 9'b000000000, 9'b111111101, 9'b111111001, 9'b000000010, 9'b000000000, 9'b000000111, 9'b000001100, 9'b111111111, 9'b000000000, 9'b000000011, 9'b111110101, 9'b111111010, 9'b000000000, 9'b000000001, 9'b111111011, 9'b000000011, 9'b000000010, 9'b111111101, 9'b111111001, 9'b111111111, 9'b000000000, 9'b111111101, 9'b000000000, 9'b000000011, 9'b111111110, 9'b000000000, 9'b000000000, 9'b111111100, 9'b111111001, 9'b000000110, 9'b000000010, 9'b111111101, 9'b000000010, 9'b111111111, 9'b111111000, 9'b111111101, 9'b111111111, 9'b111111110, 9'b000001101, 9'b000000011, 9'b111111111, 9'b111111111}, 
{9'b000000000, 9'b000001001, 9'b111110110, 9'b111111100, 9'b000000101, 9'b111111100, 9'b000010011, 9'b111111011, 9'b111111111, 9'b000000100, 9'b000000100, 9'b111111111, 9'b111111111, 9'b111111000, 9'b000000100, 9'b000000010, 9'b111111100, 9'b111111111, 9'b000000000, 9'b000000000, 9'b000000100, 9'b111111000, 9'b000000110, 9'b000001001, 9'b111111110, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000001011, 9'b000000000, 9'b111111011, 9'b000000000, 9'b000000110, 9'b111110011, 9'b111110111, 9'b000000011, 9'b000000010, 9'b111110110, 9'b111111100, 9'b111111100, 9'b000000110, 9'b000000110, 9'b000000000, 9'b111111011, 9'b000000000, 9'b000000110, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000011, 9'b111111111, 9'b111111100, 9'b000000101, 9'b111111100, 9'b000000100, 9'b000001001, 9'b000000000, 9'b000000100, 9'b111111001, 9'b111111010, 9'b000001101, 9'b111111101, 9'b000000000, 9'b111111110}, 
{9'b000000000, 9'b111111000, 9'b000000101, 9'b111111011, 9'b111111111, 9'b000000011, 9'b111110110, 9'b000000011, 9'b000000111, 9'b000000010, 9'b000000101, 9'b000000101, 9'b111111011, 9'b111111110, 9'b111111111, 9'b000000000, 9'b111110000, 9'b000000101, 9'b111111111, 9'b000000000, 9'b111111010, 9'b000000001, 9'b000000010, 9'b111111111, 9'b111111000, 9'b111111111, 9'b111111110, 9'b000010011, 9'b111110101, 9'b000000001, 9'b000000001, 9'b111111111, 9'b111111100, 9'b000000001, 9'b111111110, 9'b111111101, 9'b111111101, 9'b111111100, 9'b111111111, 9'b111111011, 9'b000000101, 9'b000000001, 9'b000000111, 9'b000000001, 9'b000000000, 9'b111111011, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000011, 9'b000000010, 9'b000000100, 9'b111111111, 9'b111111011, 9'b000000000, 9'b000000000, 9'b000000101, 9'b111111100, 9'b111110111, 9'b000001000, 9'b111111011, 9'b000010010, 9'b111111111, 9'b111111010}, 
{9'b111110110, 9'b111111111, 9'b111111001, 9'b000000011, 9'b000000100, 9'b111111110, 9'b000001000, 9'b111111101, 9'b111111000, 9'b111111010, 9'b111111011, 9'b111111000, 9'b111111100, 9'b000000011, 9'b000000000, 9'b000000000, 9'b000001101, 9'b111111111, 9'b111111111, 9'b000000110, 9'b000000100, 9'b111110110, 9'b111111001, 9'b000000011, 9'b111111001, 9'b111111111, 9'b111111011, 9'b111111010, 9'b111111001, 9'b000000100, 9'b000000011, 9'b111111101, 9'b111111110, 9'b111110000, 9'b111111101, 9'b000000000, 9'b111111101, 9'b111111011, 9'b111111111, 9'b000000001, 9'b111111110, 9'b111111111, 9'b111111111, 9'b111110101, 9'b000000000, 9'b000000000, 9'b000000101, 9'b111111110, 9'b000000110, 9'b111111100, 9'b000000100, 9'b111111111, 9'b000000011, 9'b111111001, 9'b111111111, 9'b000001000, 9'b000000101, 9'b000000100, 9'b000000000, 9'b111111001, 9'b111111011, 9'b111110101, 9'b111111111, 9'b000000001}, 
{9'b000000100, 9'b000000000, 9'b000000010, 9'b111111111, 9'b000000010, 9'b111111101, 9'b000000011, 9'b000000000, 9'b000000010, 9'b000000101, 9'b111111011, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111110101, 9'b111111011, 9'b000001010, 9'b111111111, 9'b111111111, 9'b000000000, 9'b111111001, 9'b000000000, 9'b000000100, 9'b000000000, 9'b000000000, 9'b000000101, 9'b000000000, 9'b000000000, 9'b000000000, 9'b111111111, 9'b111111100, 9'b111110101, 9'b000000100, 9'b000000101, 9'b111111111, 9'b111111100, 9'b000000000, 9'b111110101, 9'b111111111, 9'b111111111, 9'b000000011, 9'b111111101, 9'b111111111, 9'b000001101, 9'b000000111, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111100, 9'b000000010, 9'b000000010, 9'b000000010, 9'b000000010, 9'b000000110, 9'b000000101, 9'b000001010, 9'b111111101, 9'b000000110, 9'b000000010, 9'b111111010, 9'b000000001, 9'b111111001, 9'b111111000, 9'b111111000}, 
{9'b000000000, 9'b000000011, 9'b111111100, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111110101, 9'b111111111, 9'b000000100, 9'b000000011, 9'b000000011, 9'b111111001, 9'b111111110, 9'b000000100, 9'b111111111, 9'b000000000, 9'b111110010, 9'b111111111, 9'b000000101, 9'b000000001, 9'b000000011, 9'b111111110, 9'b000000011, 9'b000000110, 9'b111111010, 9'b111111011, 9'b111111111, 9'b111111110, 9'b000000001, 9'b000000000, 9'b111111111, 9'b000000101, 9'b111110100, 9'b000000101, 9'b000001000, 9'b000000001, 9'b000000001, 9'b111111110, 9'b000000001, 9'b111111110, 9'b111111011, 9'b111111111, 9'b000000010, 9'b000001011, 9'b111110010, 9'b111111000, 9'b000000011, 9'b111111110, 9'b000000111, 9'b111111100, 9'b111111010, 9'b111111011, 9'b111111111, 9'b000000001, 9'b111111101, 9'b111110010, 9'b111111101, 9'b111111111, 9'b000000000, 9'b111110110, 9'b000010001, 9'b111110111, 9'b000001000, 9'b000000010}, 
{9'b000000001, 9'b111111100, 9'b000001010, 9'b111111011, 9'b111111000, 9'b000000001, 9'b000000100, 9'b000000100, 9'b111111101, 9'b111111101, 9'b000000000, 9'b000000011, 9'b000000011, 9'b000000000, 9'b111111100, 9'b000000010, 9'b000000111, 9'b111111111, 9'b111111011, 9'b000000000, 9'b000000001, 9'b000000000, 9'b111111011, 9'b000000001, 9'b000001100, 9'b000000000, 9'b000000010, 9'b111110011, 9'b111111110, 9'b000000000, 9'b111111100, 9'b111111011, 9'b000000111, 9'b111111111, 9'b111111111, 9'b111111011, 9'b000000010, 9'b000000100, 9'b111111111, 9'b111111111, 9'b111111101, 9'b000000011, 9'b000000000, 9'b111110101, 9'b000000100, 9'b000000110, 9'b111111111, 9'b000000000, 9'b111111001, 9'b111111110, 9'b111111111, 9'b111111010, 9'b000000000, 9'b111111101, 9'b000000000, 9'b111110010, 9'b111111111, 9'b111111111, 9'b000000100, 9'b000001001, 9'b111110100, 9'b000001000, 9'b000000000, 9'b111111110}, 
{9'b000000100, 9'b000010011, 9'b000000111, 9'b000000100, 9'b111111000, 9'b111111010, 9'b111010110, 9'b111111000, 9'b000000110, 9'b111111111, 9'b000000100, 9'b000001101, 9'b000000001, 9'b000000000, 9'b111111111, 9'b000000000, 9'b111111100, 9'b111111100, 9'b000000011, 9'b111110111, 9'b111110101, 9'b111111110, 9'b111110110, 9'b000000000, 9'b111011011, 9'b000001101, 9'b000001111, 9'b000001001, 9'b111100100, 9'b111111010, 9'b111110100, 9'b111110010, 9'b111010111, 9'b000001010, 9'b111111111, 9'b000000101, 9'b000000000, 9'b111101001, 9'b000000000, 9'b000000000, 9'b000000000, 9'b000010000, 9'b111111100, 9'b111110101, 9'b000001110, 9'b111111000, 9'b111111010, 9'b111111001, 9'b000000111, 9'b000001000, 9'b111111110, 9'b111111010, 9'b111111111, 9'b111111110, 9'b000000000, 9'b111111001, 9'b000001001, 9'b000010001, 9'b000001011, 9'b111110001, 9'b111000100, 9'b000001110, 9'b000000001, 9'b000000101}, 
{9'b111111100, 9'b000000101, 9'b000000101, 9'b111111111, 9'b111111010, 9'b111111110, 9'b111111001, 9'b111111111, 9'b000000010, 9'b111111110, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111101, 9'b111111111, 9'b111111110, 9'b000000101, 9'b111111111, 9'b111110101, 9'b000000111, 9'b000001001, 9'b000000110, 9'b111111010, 9'b111111101, 9'b111111010, 9'b111111011, 9'b000000011, 9'b000000011, 9'b000000011, 9'b000000101, 9'b000000000, 9'b000000110, 9'b111111111, 9'b000000000, 9'b000000100, 9'b000000010, 9'b111111110, 9'b111111111, 9'b000000000, 9'b111111011, 9'b111111100, 9'b111111110, 9'b111111010, 9'b000000111, 9'b000000000, 9'b111111111, 9'b111111110, 9'b111111101, 9'b111110011, 9'b111111111, 9'b111111100, 9'b111111101, 9'b111111110, 9'b000000100, 9'b000001010, 9'b000000010, 9'b111111111, 9'b111111010, 9'b111111111, 9'b000000000, 9'b000000101, 9'b111111111, 9'b000000000, 9'b000000000}
};

localparam logic signed [8:0] bias [64] = '{
9'b111111111,  // -0.037350185215473175
9'b000000100,  // 0.27355897426605225
9'b111111110,  // -0.12378914654254913
9'b111111110,  // -0.064457006752491
9'b000000000,  // 0.05452875792980194
9'b000000001,  // 0.11671770364046097
9'b000000010,  // 0.13640816509723663
9'b000000001,  // 0.07482525706291199
9'b000000000,  // 0.04674031585454941
9'b111111100,  // -0.20146161317825317
9'b111111110,  // -0.09910125285387039
9'b000000010,  // 0.15104414522647858
9'b111111110,  // -0.10221704095602036
9'b111111101,  // -0.1461549550294876
9'b111111110,  // -0.08641516417264938
9'b000000010,  // 0.16613510251045227
9'b111111110,  // -0.0836295336484909
9'b111111111,  // -0.05756539851427078
9'b111111111,  // -0.03229188174009323
9'b111111111,  // -0.028388574719429016
9'b000000010,  // 0.1260243058204651
9'b111111111,  // -0.037064336240291595
9'b000000011,  // 0.19336333870887756
9'b000000000,  // 0.02124214917421341
9'b000000111,  // 0.4985624849796295
9'b000000000,  // 0.0158411655575037
9'b111111110,  // -0.08296407759189606
9'b000000001,  // 0.11056788265705109
9'b000000000,  // 0.01173810102045536
9'b111111110,  // -0.10843746364116669
9'b000000100,  // 0.27439257502555847
9'b000000001,  // 0.09199801832437515
9'b000000100,  // 0.27419957518577576
9'b000000100,  // 0.27063727378845215
9'b111111100,  // -0.24828937649726868
9'b000000001,  // 0.07818280160427094
9'b111111111,  // -0.005749030504375696
9'b000000001,  // 0.10850494354963303
9'b000000010,  // 0.13591453433036804
9'b111111110,  // -0.12088628858327866
9'b111111111,  // -0.05666546896100044
9'b000000001,  // 0.09311636537313461
9'b000000000,  // 0.05477767437696457
9'b000000000,  // 0.029585206881165504
9'b111111011,  // -0.31209176778793335
9'b111111110,  // -0.08465463668107986
9'b111111101,  // -0.16775836050510406
9'b000000010,  // 0.14762157201766968
9'b111111100,  // -0.23618532717227936
9'b000000001,  // 0.06535740196704865
9'b111111101,  // -0.12853026390075684
9'b111111101,  // -0.13802281022071838
9'b111111101,  // -0.15156887471675873
9'b000000001,  // 0.07979883998632431
9'b000000010,  // 0.18141601979732513
9'b111111111,  // -0.054039113223552704
9'b111111111,  // -0.010052933357656002
9'b000000001,  // 0.06611225008964539
9'b000000000,  // 0.05053366720676422
9'b000000000,  // 0.026860840618610382
9'b000000000,  // 0.03283466026186943
9'b000000010,  // 0.15558314323425293
9'b111111011,  // -0.2863388657569885
9'b111111110   // -0.08769102394580841
};
endpackage