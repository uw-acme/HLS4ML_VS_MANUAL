// Width: 9
// NFRAC: 4
package dense_3_9_4;

localparam logic signed [8:0] weights [32][32] = '{ 
{9'b111111111, 9'b111111001, 9'b111111001, 9'b111111100, 9'b000000101, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000010, 9'b111110111, 9'b111111111, 9'b000001101, 9'b111111100, 9'b111110001, 9'b111111111, 9'b000000001, 9'b000000110, 9'b111111010, 9'b111101110, 9'b111111111, 9'b000000000, 9'b111111001, 9'b000000000, 9'b000010000, 9'b111101000, 9'b111111100, 9'b111111001, 9'b111111101, 9'b000000110, 9'b111111101}, 
{9'b000001011, 9'b000011011, 9'b000000110, 9'b111110101, 9'b000000011, 9'b111111011, 9'b111111110, 9'b000010001, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111110110, 9'b111111100, 9'b000001000, 9'b111011110, 9'b111111000, 9'b111111111, 9'b111111111, 9'b111111111, 9'b111111101, 9'b111111011, 9'b111111011, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111101110, 9'b000000000, 9'b000000111, 9'b111111110, 9'b111110100, 9'b000000000, 9'b000000000}, 
{9'b111110000, 9'b000000010, 9'b000000000, 9'b000000101, 9'b111110101, 9'b000000000, 9'b000000000, 9'b111110010, 9'b000001000, 9'b111111011, 9'b111111011, 9'b111101000, 9'b111111011, 9'b000001000, 9'b000000100, 9'b111111111, 9'b111111110, 9'b111111111, 9'b111110010, 9'b000000000, 9'b000000001, 9'b000000001, 9'b000000011, 9'b000001110, 9'b000000000, 9'b111110011, 9'b000001100, 9'b000000000, 9'b000000010, 9'b111111111, 9'b000000000, 9'b000100100}, 
{9'b000001101, 9'b111111111, 9'b111111100, 9'b000010100, 9'b000010011, 9'b000000000, 9'b000000001, 9'b000001101, 9'b111111001, 9'b111111111, 9'b111110010, 9'b000000001, 9'b000000100, 9'b111110100, 9'b000000001, 9'b111111101, 9'b111111111, 9'b111111010, 9'b000000000, 9'b000000000, 9'b000000000, 9'b111111110, 9'b000010011, 9'b000001010, 9'b000001010, 9'b000000111, 9'b000001010, 9'b000000000, 9'b111111110, 9'b000001110, 9'b000000111, 9'b111111101}, 
{9'b000010000, 9'b111111110, 9'b111110100, 9'b111100111, 9'b000001111, 9'b000000000, 9'b111110010, 9'b111110110, 9'b111111110, 9'b111100110, 9'b111011100, 9'b000001111, 9'b000010101, 9'b000010000, 9'b111101101, 9'b111100111, 9'b000000000, 9'b111111011, 9'b000000110, 9'b000000100, 9'b111111001, 9'b111111111, 9'b000010111, 9'b111010100, 9'b000000010, 9'b111101010, 9'b000000010, 9'b111111000, 9'b111110110, 9'b111111111, 9'b000000010, 9'b000010010}, 
{9'b000000001, 9'b111111110, 9'b111110110, 9'b111110111, 9'b000001011, 9'b000000000, 9'b111110111, 9'b111111011, 9'b111110010, 9'b111111101, 9'b111111111, 9'b000000101, 9'b000000000, 9'b000001011, 9'b111101111, 9'b111111011, 9'b000000010, 9'b111110110, 9'b111111001, 9'b111111111, 9'b000000000, 9'b000001001, 9'b000001110, 9'b111111111, 9'b111111111, 9'b000001100, 9'b111101110, 9'b111111111, 9'b111111000, 9'b111111110, 9'b111111111, 9'b000000000}, 
{9'b000000010, 9'b111110101, 9'b000000011, 9'b111111110, 9'b111111111, 9'b000000100, 9'b111111100, 9'b111101010, 9'b111111111, 9'b111111001, 9'b111110001, 9'b000001111, 9'b000000000, 9'b000010101, 9'b000011010, 9'b000000000, 9'b111111111, 9'b111110101, 9'b111111110, 9'b000001000, 9'b111100111, 9'b000000100, 9'b000001010, 9'b000000000, 9'b000000100, 9'b000100111, 9'b111110011, 9'b111111101, 9'b111111001, 9'b000001111, 9'b111111110, 9'b111111010}, 
{9'b111101100, 9'b000000000, 9'b111101011, 9'b000001101, 9'b000100000, 9'b000000011, 9'b000000000, 9'b000000001, 9'b111111111, 9'b000000100, 9'b000101001, 9'b111111111, 9'b000001100, 9'b000010011, 9'b000011000, 9'b000100001, 9'b000000000, 9'b111110000, 9'b000001010, 9'b111111111, 9'b111101011, 9'b111111000, 9'b000000000, 9'b111111101, 9'b111101111, 9'b000111100, 9'b111111000, 9'b000000000, 9'b000000000, 9'b000011100, 9'b000000010, 9'b000001100}, 
{9'b000001101, 9'b111111111, 9'b000000000, 9'b111111110, 9'b000000010, 9'b111111110, 9'b111111111, 9'b000000101, 9'b000000110, 9'b111110111, 9'b000000100, 9'b000000101, 9'b000000000, 9'b000001010, 9'b111111000, 9'b111100110, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111110000, 9'b111111111, 9'b000000000, 9'b111111001, 9'b111111111, 9'b111111100, 9'b000000100, 9'b000001011, 9'b111111100, 9'b111111110, 9'b111111110, 9'b000000000, 9'b111110011}, 
{9'b111111010, 9'b000001100, 9'b000000000, 9'b000000000, 9'b000011001, 9'b000001010, 9'b111111111, 9'b111101110, 9'b000000011, 9'b111101001, 9'b111010011, 9'b111111111, 9'b000000000, 9'b000001101, 9'b000000011, 9'b000000000, 9'b111110101, 9'b000000000, 9'b000000000, 9'b000000001, 9'b000000111, 9'b111111111, 9'b111110100, 9'b000000000, 9'b111111111, 9'b000100010, 9'b000001010, 9'b111111111, 9'b111111101, 9'b000010101, 9'b111111110, 9'b111111101}, 
{9'b111101111, 9'b000000101, 9'b111111110, 9'b111111111, 9'b111111000, 9'b111110011, 9'b000000001, 9'b000000100, 9'b111111111, 9'b111111010, 9'b111101101, 9'b000000110, 9'b000001001, 9'b000000000, 9'b000011010, 9'b111101110, 9'b000000011, 9'b111110011, 9'b000001001, 9'b111111111, 9'b111111110, 9'b000000010, 9'b000000011, 9'b000000000, 9'b111110000, 9'b000000000, 9'b111101110, 9'b111111110, 9'b111111111, 9'b000010101, 9'b111111001, 9'b000000000}, 
{9'b111111111, 9'b000000011, 9'b000000000, 9'b000001100, 9'b111111100, 9'b111111110, 9'b000000001, 9'b111111111, 9'b111111110, 9'b000010100, 9'b000010110, 9'b000000000, 9'b111110101, 9'b111101001, 9'b111111110, 9'b000000000, 9'b000000000, 9'b111111101, 9'b111110000, 9'b000001100, 9'b000000000, 9'b000001011, 9'b111111111, 9'b000010001, 9'b000000011, 9'b000001001, 9'b000001110, 9'b111111110, 9'b111110011, 9'b111110001, 9'b111111111, 9'b111101010}, 
{9'b111111000, 9'b111111111, 9'b000000011, 9'b111110010, 9'b000000010, 9'b111111111, 9'b111111001, 9'b111111111, 9'b111111011, 9'b000000001, 9'b000000010, 9'b111111101, 9'b000000000, 9'b000000110, 9'b111101011, 9'b111111000, 9'b000000111, 9'b111111010, 9'b000000000, 9'b111111111, 9'b000000110, 9'b000000000, 9'b111111111, 9'b000000001, 9'b000001000, 9'b111111100, 9'b000000000, 9'b111110001, 9'b111111001, 9'b111111111, 9'b000000101, 9'b000000000}, 
{9'b111101111, 9'b000001101, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000101, 9'b111111111, 9'b000011000, 9'b111111111, 9'b111111111, 9'b000000110, 9'b000000001, 9'b000000000, 9'b000000000, 9'b000000011, 9'b000001010, 9'b000000101, 9'b000000101, 9'b111111111, 9'b000001001, 9'b000000011, 9'b000000001, 9'b111111111, 9'b000001000, 9'b111111100, 9'b111110101, 9'b111111101, 9'b111111111, 9'b000000011, 9'b000000000, 9'b000000110, 9'b000001111}, 
{9'b111111111, 9'b111110011, 9'b000000001, 9'b111111111, 9'b000011101, 9'b111111001, 9'b111101101, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000001, 9'b000001101, 9'b000001010, 9'b000000000, 9'b000000001, 9'b111111010, 9'b000000001, 9'b111111110, 9'b000000000, 9'b000000010, 9'b111111110, 9'b000000000, 9'b000001000, 9'b000000001, 9'b111111111, 9'b111110010, 9'b000000110, 9'b111111111, 9'b111111111, 9'b111111100, 9'b111111111, 9'b111111101}, 
{9'b000000000, 9'b111111101, 9'b111111011, 9'b111111001, 9'b111101110, 9'b000010011, 9'b000000000, 9'b000000101, 9'b000001001, 9'b000000000, 9'b111111110, 9'b000001111, 9'b000000111, 9'b111110100, 9'b111111010, 9'b111111110, 9'b111110011, 9'b111111111, 9'b000000000, 9'b111111111, 9'b000000100, 9'b111111011, 9'b000000000, 9'b000000010, 9'b111111111, 9'b111110101, 9'b000000101, 9'b000000000, 9'b000000001, 9'b000000000, 9'b111110101, 9'b000000000}, 
{9'b111111001, 9'b111111010, 9'b000000010, 9'b111111100, 9'b111111101, 9'b000000011, 9'b111111111, 9'b000000001, 9'b000000100, 9'b111111111, 9'b000000011, 9'b111111011, 9'b111111111, 9'b111111111, 9'b000000011, 9'b111111111, 9'b000001111, 9'b111111111, 9'b000000111, 9'b111111010, 9'b000000101, 9'b000000010, 9'b000000010, 9'b000000001, 9'b111111101, 9'b111110111, 9'b111110111, 9'b000000011, 9'b111111101, 9'b000000000, 9'b111111111, 9'b000000111}, 
{9'b111111111, 9'b111110011, 9'b111110011, 9'b111111111, 9'b000010100, 9'b111111101, 9'b000000000, 9'b000001111, 9'b111111011, 9'b000000000, 9'b111110010, 9'b111110000, 9'b000001110, 9'b000000100, 9'b111111100, 9'b111110111, 9'b000000101, 9'b000000000, 9'b111111000, 9'b000000000, 9'b000000010, 9'b111111101, 9'b000001001, 9'b111100000, 9'b000000001, 9'b000000111, 9'b111111110, 9'b000000000, 9'b111111000, 9'b111111111, 9'b111111001, 9'b111111111}, 
{9'b000000110, 9'b000001011, 9'b000010001, 9'b111111001, 9'b000001101, 9'b000001001, 9'b000000000, 9'b000001110, 9'b000001011, 9'b111111100, 9'b000010110, 9'b111110100, 9'b000010011, 9'b000001110, 9'b111011101, 9'b111111111, 9'b000000000, 9'b000000000, 9'b000001000, 9'b111101111, 9'b000000111, 9'b111111001, 9'b111110000, 9'b111111010, 9'b000001010, 9'b111101010, 9'b111110101, 9'b111111110, 9'b111111111, 9'b111101101, 9'b000001100, 9'b000000000}, 
{9'b111111110, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111110100, 9'b000000000, 9'b000000000, 9'b111111111, 9'b111111111, 9'b111111110, 9'b000000100, 9'b111111111, 9'b000000010, 9'b111110101, 9'b000000011, 9'b111111111, 9'b000000100, 9'b000001110, 9'b111110100, 9'b000000001, 9'b111111100, 9'b000000100, 9'b000000110, 9'b111111101, 9'b111110111, 9'b000000000, 9'b000011010, 9'b111111111, 9'b111111111, 9'b000001010, 9'b000000000, 9'b000011011}, 
{9'b111101111, 9'b000000001, 9'b111111001, 9'b000001100, 9'b000000011, 9'b111111110, 9'b111111111, 9'b111111111, 9'b111110110, 9'b111111110, 9'b000000000, 9'b111101110, 9'b000000000, 9'b111111110, 9'b111111111, 9'b111111111, 9'b111111100, 9'b000000000, 9'b000000000, 9'b000000101, 9'b000000000, 9'b000000000, 9'b000000000, 9'b111111111, 9'b000000000, 9'b000000000, 9'b000010010, 9'b111111111, 9'b111111111, 9'b111111110, 9'b000000101, 9'b111111111}, 
{9'b111111111, 9'b111111011, 9'b000000110, 9'b000000001, 9'b111110100, 9'b000000000, 9'b000001001, 9'b111111111, 9'b000000000, 9'b111111100, 9'b000000011, 9'b000000000, 9'b000001010, 9'b111101110, 9'b111111100, 9'b111111111, 9'b000000110, 9'b111110011, 9'b000000000, 9'b111100111, 9'b111111111, 9'b111111100, 9'b111111110, 9'b000001001, 9'b111111101, 9'b111110111, 9'b000000010, 9'b000000000, 9'b000001100, 9'b000010000, 9'b111110101, 9'b111110001}, 
{9'b000000010, 9'b000000000, 9'b111110010, 9'b111111110, 9'b111111111, 9'b000000000, 9'b000000011, 9'b000001101, 9'b000000000, 9'b000000000, 9'b000000010, 9'b111101110, 9'b111111101, 9'b111101100, 9'b000001111, 9'b000000000, 9'b111111111, 9'b111101011, 9'b111111111, 9'b111111101, 9'b111111111, 9'b000000000, 9'b000000001, 9'b111111011, 9'b000000001, 9'b000001101, 9'b000001101, 9'b000001100, 9'b000001001, 9'b000000000, 9'b000000011, 9'b000011001}, 
{9'b111111111, 9'b111111000, 9'b000001100, 9'b111111100, 9'b000000010, 9'b000000101, 9'b111111111, 9'b111110110, 9'b111111101, 9'b111101100, 9'b000001110, 9'b000000000, 9'b000001101, 9'b000010101, 9'b111111100, 9'b111100100, 9'b111111100, 9'b000001111, 9'b111110110, 9'b111111001, 9'b000000001, 9'b000000000, 9'b111101110, 9'b111111001, 9'b111111110, 9'b111111100, 9'b000000011, 9'b000010110, 9'b000000111, 9'b111111111, 9'b000000010, 9'b000000000}, 
{9'b000000001, 9'b000001110, 9'b000000000, 9'b000001001, 9'b000011010, 9'b111111010, 9'b111111111, 9'b111111110, 9'b000001001, 9'b111111001, 9'b111111111, 9'b000001010, 9'b000000000, 9'b000000000, 9'b111001111, 9'b111111101, 9'b000000000, 9'b000000110, 9'b111111111, 9'b000001001, 9'b111111111, 9'b111111010, 9'b111101110, 9'b000000100, 9'b000001001, 9'b111011100, 9'b111111111, 9'b000000000, 9'b000010001, 9'b111100110, 9'b000000000, 9'b111111111}, 
{9'b000000000, 9'b111110101, 9'b000000001, 9'b111111111, 9'b000000001, 9'b000010000, 9'b111101000, 9'b000000001, 9'b000001101, 9'b111110101, 9'b111111111, 9'b000000001, 9'b111111111, 9'b000000101, 9'b000000011, 9'b111111111, 9'b000000010, 9'b000000000, 9'b000000000, 9'b000001100, 9'b111111111, 9'b111110000, 9'b111101100, 9'b111111001, 9'b111101101, 9'b000000110, 9'b000010011, 9'b000001011, 9'b111111111, 9'b111110100, 9'b111110110, 9'b000000001}, 
{9'b000000001, 9'b111110000, 9'b111111111, 9'b000000100, 9'b111110000, 9'b000000101, 9'b111111111, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000001000, 9'b111111111, 9'b000000000, 9'b000000000, 9'b000000100, 9'b111111111, 9'b000000000, 9'b111111111, 9'b111110101, 9'b111101111, 9'b111111111, 9'b111101110, 9'b111110110, 9'b111110100, 9'b000011100, 9'b000000000, 9'b111111110, 9'b000001010, 9'b000011100, 9'b000001100, 9'b111011110, 9'b111111010}, 
{9'b000001100, 9'b111111111, 9'b000001000, 9'b111111111, 9'b000001111, 9'b111111011, 9'b000000010, 9'b000001101, 9'b000001000, 9'b111101111, 9'b111111110, 9'b000000011, 9'b000000010, 9'b111111111, 9'b000000010, 9'b000000000, 9'b000001011, 9'b000000001, 9'b000001011, 9'b111111101, 9'b111111011, 9'b111111101, 9'b111111111, 9'b000001001, 9'b111111001, 9'b111111111, 9'b000000000, 9'b000000000, 9'b000000000, 9'b000001001, 9'b111110101, 9'b111111111}, 
{9'b111111111, 9'b111111111, 9'b111110001, 9'b000001001, 9'b000000111, 9'b111111100, 9'b111111111, 9'b111111000, 9'b000000000, 9'b111111111, 9'b111110110, 9'b111111000, 9'b000001111, 9'b000000000, 9'b111111011, 9'b111111111, 9'b000000110, 9'b111111111, 9'b111111111, 9'b111111001, 9'b000001010, 9'b000000000, 9'b000000100, 9'b111111111, 9'b000000101, 9'b000000000, 9'b000000000, 9'b000000111, 9'b111111001, 9'b111111110, 9'b000000101, 9'b111111100}, 
{9'b111111111, 9'b111110110, 9'b000010011, 9'b111111101, 9'b000000110, 9'b111110110, 9'b000000000, 9'b000000001, 9'b111110000, 9'b111111111, 9'b111111100, 9'b000000001, 9'b111110101, 9'b000000100, 9'b000000110, 9'b000000011, 9'b000000010, 9'b111111110, 9'b111101001, 9'b111111111, 9'b111111110, 9'b000000100, 9'b111111100, 9'b111111111, 9'b000000110, 9'b111111110, 9'b111111111, 9'b000001100, 9'b111110011, 9'b111110110, 9'b000001011, 9'b000000001}, 
{9'b000001101, 9'b000000110, 9'b000000000, 9'b111111010, 9'b111111101, 9'b111111111, 9'b000000000, 9'b111111101, 9'b111111100, 9'b111111100, 9'b000000000, 9'b000000101, 9'b000000000, 9'b000000001, 9'b111111110, 9'b000000000, 9'b111111011, 9'b000000000, 9'b111111111, 9'b111111111, 9'b000000000, 9'b000000001, 9'b000000011, 9'b000000000, 9'b000000000, 9'b111101100, 9'b111111001, 9'b000000000, 9'b000000000, 9'b000000000, 9'b111111010, 9'b000000000}, 
{9'b000000110, 9'b111011110, 9'b111111111, 9'b111111101, 9'b111111000, 9'b111111111, 9'b000000000, 9'b000010001, 9'b111111110, 9'b111111111, 9'b000000010, 9'b111101010, 9'b000000000, 9'b111110001, 9'b000010111, 9'b111111110, 9'b111111000, 9'b111101110, 9'b111111111, 9'b111101001, 9'b111100110, 9'b111111111, 9'b000000000, 9'b000000000, 9'b000000111, 9'b111111111, 9'b111110110, 9'b111111101, 9'b111111111, 9'b000000000, 9'b111111110, 9'b111101001}
};

localparam logic signed [8:0] bias [32] = '{
9'b000001000,  // 0.5280959606170654
9'b000001101,  // 0.8414360880851746
9'b000000110,  // 0.397830605506897
9'b000000110,  // 0.4105983078479767
9'b111000101,  // -3.657735586166382
9'b111110001,  // -0.8977976441383362
9'b000011011,  // 1.7051936388015747
9'b111101011,  // -1.2765135765075684
9'b111110110,  // -0.5837795734405518
9'b000101011,  // 2.699671983718872
9'b000000011,  // 0.2170683741569519
9'b000001110,  // 0.8814588785171509
9'b111010101,  // -2.634300947189331
9'b111100001,  // -1.877297282218933
9'b000011010,  // 1.6625694036483765
9'b000101011,  // 2.7459704875946045
9'b111111000,  // -0.47838035225868225
9'b000011011,  // 1.6984987258911133
9'b000001101,  // 0.8548859357833862
9'b000010000,  // 1.0045719146728516
9'b000010110,  // 1.4197649955749512
9'b000001101,  // 0.832463800907135
9'b000001000,  // 0.5434179306030273
9'b000001110,  // 0.9277304410934448
9'b111111010,  // -0.3426123857498169
9'b111110111,  // -0.5587119460105896
9'b111110110,  // -0.6208624839782715
9'b111101011,  // -1.2802538871765137
9'b000000000,  // 0.05940237268805504
9'b111110010,  // -0.8213341236114502
9'b000001110,  // 0.8783953189849854
9'b111110000   // -0.949700653553009
};
endpackage