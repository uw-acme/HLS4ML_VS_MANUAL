// Width: 8
// NFRAC: 4
package dense_3_8_4;

localparam logic signed [7:0] weights [32][32] = '{ 
{8'b11111111, 8'b11111001, 8'b11111001, 8'b11111100, 8'b00000101, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000010, 8'b11110111, 8'b11111111, 8'b00001101, 8'b11111100, 8'b11110001, 8'b11111111, 8'b00000001, 8'b00000110, 8'b11111010, 8'b11101110, 8'b11111111, 8'b00000000, 8'b11111001, 8'b00000000, 8'b00010000, 8'b11101000, 8'b11111100, 8'b11111001, 8'b11111101, 8'b00000110, 8'b11111101}, 
{8'b00001011, 8'b00011011, 8'b00000110, 8'b11110101, 8'b00000011, 8'b11111011, 8'b11111110, 8'b00010001, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11110110, 8'b11111100, 8'b00001000, 8'b11011110, 8'b11111000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111101, 8'b11111011, 8'b11111011, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11101110, 8'b00000000, 8'b00000111, 8'b11111110, 8'b11110100, 8'b00000000, 8'b00000000}, 
{8'b11110000, 8'b00000010, 8'b00000000, 8'b00000101, 8'b11110101, 8'b00000000, 8'b00000000, 8'b11110010, 8'b00001000, 8'b11111011, 8'b11111011, 8'b11101000, 8'b11111011, 8'b00001000, 8'b00000100, 8'b11111111, 8'b11111110, 8'b11111111, 8'b11110010, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000011, 8'b00001110, 8'b00000000, 8'b11110011, 8'b00001100, 8'b00000000, 8'b00000010, 8'b11111111, 8'b00000000, 8'b00100100}, 
{8'b00001101, 8'b11111111, 8'b11111100, 8'b00010100, 8'b00010011, 8'b00000000, 8'b00000001, 8'b00001101, 8'b11111001, 8'b11111111, 8'b11110010, 8'b00000001, 8'b00000100, 8'b11110100, 8'b00000001, 8'b11111101, 8'b11111111, 8'b11111010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111110, 8'b00010011, 8'b00001010, 8'b00001010, 8'b00000111, 8'b00001010, 8'b00000000, 8'b11111110, 8'b00001110, 8'b00000111, 8'b11111101}, 
{8'b00010000, 8'b11111110, 8'b11110100, 8'b11100111, 8'b00001111, 8'b00000000, 8'b11110010, 8'b11110110, 8'b11111110, 8'b11100110, 8'b11011100, 8'b00001111, 8'b00010101, 8'b00010000, 8'b11101101, 8'b11100111, 8'b00000000, 8'b11111011, 8'b00000110, 8'b00000100, 8'b11111001, 8'b11111111, 8'b00010111, 8'b11010100, 8'b00000010, 8'b11101010, 8'b00000010, 8'b11111000, 8'b11110110, 8'b11111111, 8'b00000010, 8'b00010010}, 
{8'b00000001, 8'b11111110, 8'b11110110, 8'b11110111, 8'b00001011, 8'b00000000, 8'b11110111, 8'b11111011, 8'b11110010, 8'b11111101, 8'b11111111, 8'b00000101, 8'b00000000, 8'b00001011, 8'b11101111, 8'b11111011, 8'b00000010, 8'b11110110, 8'b11111001, 8'b11111111, 8'b00000000, 8'b00001001, 8'b00001110, 8'b11111111, 8'b11111111, 8'b00001100, 8'b11101110, 8'b11111111, 8'b11111000, 8'b11111110, 8'b11111111, 8'b00000000}, 
{8'b00000010, 8'b11110101, 8'b00000011, 8'b11111110, 8'b11111111, 8'b00000100, 8'b11111100, 8'b11101010, 8'b11111111, 8'b11111001, 8'b11110001, 8'b00001111, 8'b00000000, 8'b00010101, 8'b00011010, 8'b00000000, 8'b11111111, 8'b11110101, 8'b11111110, 8'b00001000, 8'b11100111, 8'b00000100, 8'b00001010, 8'b00000000, 8'b00000100, 8'b00100111, 8'b11110011, 8'b11111101, 8'b11111001, 8'b00001111, 8'b11111110, 8'b11111010}, 
{8'b11101100, 8'b00000000, 8'b11101011, 8'b00001101, 8'b00100000, 8'b00000011, 8'b00000000, 8'b00000001, 8'b11111111, 8'b00000100, 8'b00101001, 8'b11111111, 8'b00001100, 8'b00010011, 8'b00011000, 8'b00100001, 8'b00000000, 8'b11110000, 8'b00001010, 8'b11111111, 8'b11101011, 8'b11111000, 8'b00000000, 8'b11111101, 8'b11101111, 8'b00111100, 8'b11111000, 8'b00000000, 8'b00000000, 8'b00011100, 8'b00000010, 8'b00001100}, 
{8'b00001101, 8'b11111111, 8'b00000000, 8'b11111110, 8'b00000010, 8'b11111110, 8'b11111111, 8'b00000101, 8'b00000110, 8'b11110111, 8'b00000100, 8'b00000101, 8'b00000000, 8'b00001010, 8'b11111000, 8'b11100110, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11110000, 8'b11111111, 8'b00000000, 8'b11111001, 8'b11111111, 8'b11111100, 8'b00000100, 8'b00001011, 8'b11111100, 8'b11111110, 8'b11111110, 8'b00000000, 8'b11110011}, 
{8'b11111010, 8'b00001100, 8'b00000000, 8'b00000000, 8'b00011001, 8'b00001010, 8'b11111111, 8'b11101110, 8'b00000011, 8'b11101001, 8'b11010011, 8'b11111111, 8'b00000000, 8'b00001101, 8'b00000011, 8'b00000000, 8'b11110101, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000111, 8'b11111111, 8'b11110100, 8'b00000000, 8'b11111111, 8'b00100010, 8'b00001010, 8'b11111111, 8'b11111101, 8'b00010101, 8'b11111110, 8'b11111101}, 
{8'b11101111, 8'b00000101, 8'b11111110, 8'b11111111, 8'b11111000, 8'b11110011, 8'b00000001, 8'b00000100, 8'b11111111, 8'b11111010, 8'b11101101, 8'b00000110, 8'b00001001, 8'b00000000, 8'b00011010, 8'b11101110, 8'b00000011, 8'b11110011, 8'b00001001, 8'b11111111, 8'b11111110, 8'b00000010, 8'b00000011, 8'b00000000, 8'b11110000, 8'b00000000, 8'b11101110, 8'b11111110, 8'b11111111, 8'b00010101, 8'b11111001, 8'b00000000}, 
{8'b11111111, 8'b00000011, 8'b00000000, 8'b00001100, 8'b11111100, 8'b11111110, 8'b00000001, 8'b11111111, 8'b11111110, 8'b00010100, 8'b00010110, 8'b00000000, 8'b11110101, 8'b11101001, 8'b11111110, 8'b00000000, 8'b00000000, 8'b11111101, 8'b11110000, 8'b00001100, 8'b00000000, 8'b00001011, 8'b11111111, 8'b00010001, 8'b00000011, 8'b00001001, 8'b00001110, 8'b11111110, 8'b11110011, 8'b11110001, 8'b11111111, 8'b11101010}, 
{8'b11111000, 8'b11111111, 8'b00000011, 8'b11110010, 8'b00000010, 8'b11111111, 8'b11111001, 8'b11111111, 8'b11111011, 8'b00000001, 8'b00000010, 8'b11111101, 8'b00000000, 8'b00000110, 8'b11101011, 8'b11111000, 8'b00000111, 8'b11111010, 8'b00000000, 8'b11111111, 8'b00000110, 8'b00000000, 8'b11111111, 8'b00000001, 8'b00001000, 8'b11111100, 8'b00000000, 8'b11110001, 8'b11111001, 8'b11111111, 8'b00000101, 8'b00000000}, 
{8'b11101111, 8'b00001101, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000101, 8'b11111111, 8'b00011000, 8'b11111111, 8'b11111111, 8'b00000110, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000011, 8'b00001010, 8'b00000101, 8'b00000101, 8'b11111111, 8'b00001001, 8'b00000011, 8'b00000001, 8'b11111111, 8'b00001000, 8'b11111100, 8'b11110101, 8'b11111101, 8'b11111111, 8'b00000011, 8'b00000000, 8'b00000110, 8'b00001111}, 
{8'b11111111, 8'b11110011, 8'b00000001, 8'b11111111, 8'b00011101, 8'b11111001, 8'b11101101, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000001, 8'b00001101, 8'b00001010, 8'b00000000, 8'b00000001, 8'b11111010, 8'b00000001, 8'b11111110, 8'b00000000, 8'b00000010, 8'b11111110, 8'b00000000, 8'b00001000, 8'b00000001, 8'b11111111, 8'b11110010, 8'b00000110, 8'b11111111, 8'b11111111, 8'b11111100, 8'b11111111, 8'b11111101}, 
{8'b00000000, 8'b11111101, 8'b11111011, 8'b11111001, 8'b11101110, 8'b00010011, 8'b00000000, 8'b00000101, 8'b00001001, 8'b00000000, 8'b11111110, 8'b00001111, 8'b00000111, 8'b11110100, 8'b11111010, 8'b11111110, 8'b11110011, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000100, 8'b11111011, 8'b00000000, 8'b00000010, 8'b11111111, 8'b11110101, 8'b00000101, 8'b00000000, 8'b00000001, 8'b00000000, 8'b11110101, 8'b00000000}, 
{8'b11111001, 8'b11111010, 8'b00000010, 8'b11111100, 8'b11111101, 8'b00000011, 8'b11111111, 8'b00000001, 8'b00000100, 8'b11111111, 8'b00000011, 8'b11111011, 8'b11111111, 8'b11111111, 8'b00000011, 8'b11111111, 8'b00001111, 8'b11111111, 8'b00000111, 8'b11111010, 8'b00000101, 8'b00000010, 8'b00000010, 8'b00000001, 8'b11111101, 8'b11110111, 8'b11110111, 8'b00000011, 8'b11111101, 8'b00000000, 8'b11111111, 8'b00000111}, 
{8'b11111111, 8'b11110011, 8'b11110011, 8'b11111111, 8'b00010100, 8'b11111101, 8'b00000000, 8'b00001111, 8'b11111011, 8'b00000000, 8'b11110010, 8'b11110000, 8'b00001110, 8'b00000100, 8'b11111100, 8'b11110111, 8'b00000101, 8'b00000000, 8'b11111000, 8'b00000000, 8'b00000010, 8'b11111101, 8'b00001001, 8'b11100000, 8'b00000001, 8'b00000111, 8'b11111110, 8'b00000000, 8'b11111000, 8'b11111111, 8'b11111001, 8'b11111111}, 
{8'b00000110, 8'b00001011, 8'b00010001, 8'b11111001, 8'b00001101, 8'b00001001, 8'b00000000, 8'b00001110, 8'b00001011, 8'b11111100, 8'b00010110, 8'b11110100, 8'b00010011, 8'b00001110, 8'b11011101, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00001000, 8'b11101111, 8'b00000111, 8'b11111001, 8'b11110000, 8'b11111010, 8'b00001010, 8'b11101010, 8'b11110101, 8'b11111110, 8'b11111111, 8'b11101101, 8'b00001100, 8'b00000000}, 
{8'b11111110, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11110100, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111110, 8'b00000100, 8'b11111111, 8'b00000010, 8'b11110101, 8'b00000011, 8'b11111111, 8'b00000100, 8'b00001110, 8'b11110100, 8'b00000001, 8'b11111100, 8'b00000100, 8'b00000110, 8'b11111101, 8'b11110111, 8'b00000000, 8'b00011010, 8'b11111111, 8'b11111111, 8'b00001010, 8'b00000000, 8'b00011011}, 
{8'b11101111, 8'b00000001, 8'b11111001, 8'b00001100, 8'b00000011, 8'b11111110, 8'b11111111, 8'b11111111, 8'b11110110, 8'b11111110, 8'b00000000, 8'b11101110, 8'b00000000, 8'b11111110, 8'b11111111, 8'b11111111, 8'b11111100, 8'b00000000, 8'b00000000, 8'b00000101, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00010010, 8'b11111111, 8'b11111111, 8'b11111110, 8'b00000101, 8'b11111111}, 
{8'b11111111, 8'b11111011, 8'b00000110, 8'b00000001, 8'b11110100, 8'b00000000, 8'b00001001, 8'b11111111, 8'b00000000, 8'b11111100, 8'b00000011, 8'b00000000, 8'b00001010, 8'b11101110, 8'b11111100, 8'b11111111, 8'b00000110, 8'b11110011, 8'b00000000, 8'b11100111, 8'b11111111, 8'b11111100, 8'b11111110, 8'b00001001, 8'b11111101, 8'b11110111, 8'b00000010, 8'b00000000, 8'b00001100, 8'b00010000, 8'b11110101, 8'b11110001}, 
{8'b00000010, 8'b00000000, 8'b11110010, 8'b11111110, 8'b11111111, 8'b00000000, 8'b00000011, 8'b00001101, 8'b00000000, 8'b00000000, 8'b00000010, 8'b11101110, 8'b11111101, 8'b11101100, 8'b00001111, 8'b00000000, 8'b11111111, 8'b11101011, 8'b11111111, 8'b11111101, 8'b11111111, 8'b00000000, 8'b00000001, 8'b11111011, 8'b00000001, 8'b00001101, 8'b00001101, 8'b00001100, 8'b00001001, 8'b00000000, 8'b00000011, 8'b00011001}, 
{8'b11111111, 8'b11111000, 8'b00001100, 8'b11111100, 8'b00000010, 8'b00000101, 8'b11111111, 8'b11110110, 8'b11111101, 8'b11101100, 8'b00001110, 8'b00000000, 8'b00001101, 8'b00010101, 8'b11111100, 8'b11100100, 8'b11111100, 8'b00001111, 8'b11110110, 8'b11111001, 8'b00000001, 8'b00000000, 8'b11101110, 8'b11111001, 8'b11111110, 8'b11111100, 8'b00000011, 8'b00010110, 8'b00000111, 8'b11111111, 8'b00000010, 8'b00000000}, 
{8'b00000001, 8'b00001110, 8'b00000000, 8'b00001001, 8'b00011010, 8'b11111010, 8'b11111111, 8'b11111110, 8'b00001001, 8'b11111001, 8'b11111111, 8'b00001010, 8'b00000000, 8'b00000000, 8'b11001111, 8'b11111101, 8'b00000000, 8'b00000110, 8'b11111111, 8'b00001001, 8'b11111111, 8'b11111010, 8'b11101110, 8'b00000100, 8'b00001001, 8'b11011100, 8'b11111111, 8'b00000000, 8'b00010001, 8'b11100110, 8'b00000000, 8'b11111111}, 
{8'b00000000, 8'b11110101, 8'b00000001, 8'b11111111, 8'b00000001, 8'b00010000, 8'b11101000, 8'b00000001, 8'b00001101, 8'b11110101, 8'b11111111, 8'b00000001, 8'b11111111, 8'b00000101, 8'b00000011, 8'b11111111, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00001100, 8'b11111111, 8'b11110000, 8'b11101100, 8'b11111001, 8'b11101101, 8'b00000110, 8'b00010011, 8'b00001011, 8'b11111111, 8'b11110100, 8'b11110110, 8'b00000001}, 
{8'b00000001, 8'b11110000, 8'b11111111, 8'b00000100, 8'b11110000, 8'b00000101, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00001000, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000100, 8'b11111111, 8'b00000000, 8'b11111111, 8'b11110101, 8'b11101111, 8'b11111111, 8'b11101110, 8'b11110110, 8'b11110100, 8'b00011100, 8'b00000000, 8'b11111110, 8'b00001010, 8'b00011100, 8'b00001100, 8'b11011110, 8'b11111010}, 
{8'b00001100, 8'b11111111, 8'b00001000, 8'b11111111, 8'b00001111, 8'b11111011, 8'b00000010, 8'b00001101, 8'b00001000, 8'b11101111, 8'b11111110, 8'b00000011, 8'b00000010, 8'b11111111, 8'b00000010, 8'b00000000, 8'b00001011, 8'b00000001, 8'b00001011, 8'b11111101, 8'b11111011, 8'b11111101, 8'b11111111, 8'b00001001, 8'b11111001, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001001, 8'b11110101, 8'b11111111}, 
{8'b11111111, 8'b11111111, 8'b11110001, 8'b00001001, 8'b00000111, 8'b11111100, 8'b11111111, 8'b11111000, 8'b00000000, 8'b11111111, 8'b11110110, 8'b11111000, 8'b00001111, 8'b00000000, 8'b11111011, 8'b11111111, 8'b00000110, 8'b11111111, 8'b11111111, 8'b11111001, 8'b00001010, 8'b00000000, 8'b00000100, 8'b11111111, 8'b00000101, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11111001, 8'b11111110, 8'b00000101, 8'b11111100}, 
{8'b11111111, 8'b11110110, 8'b00010011, 8'b11111101, 8'b00000110, 8'b11110110, 8'b00000000, 8'b00000001, 8'b11110000, 8'b11111111, 8'b11111100, 8'b00000001, 8'b11110101, 8'b00000100, 8'b00000110, 8'b00000011, 8'b00000010, 8'b11111110, 8'b11101001, 8'b11111111, 8'b11111110, 8'b00000100, 8'b11111100, 8'b11111111, 8'b00000110, 8'b11111110, 8'b11111111, 8'b00001100, 8'b11110011, 8'b11110110, 8'b00001011, 8'b00000001}, 
{8'b00001101, 8'b00000110, 8'b00000000, 8'b11111010, 8'b11111101, 8'b11111111, 8'b00000000, 8'b11111101, 8'b11111100, 8'b11111100, 8'b00000000, 8'b00000101, 8'b00000000, 8'b00000001, 8'b11111110, 8'b00000000, 8'b11111011, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000001, 8'b00000011, 8'b00000000, 8'b00000000, 8'b11101100, 8'b11111001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111010, 8'b00000000}, 
{8'b00000110, 8'b11011110, 8'b11111111, 8'b11111101, 8'b11111000, 8'b11111111, 8'b00000000, 8'b00010001, 8'b11111110, 8'b11111111, 8'b00000010, 8'b11101010, 8'b00000000, 8'b11110001, 8'b00010111, 8'b11111110, 8'b11111000, 8'b11101110, 8'b11111111, 8'b11101001, 8'b11100110, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11111111, 8'b11110110, 8'b11111101, 8'b11111111, 8'b00000000, 8'b11111110, 8'b11101001}
};

localparam logic signed [7:0] bias [32] = '{
8'b00001000,  // 0.5280959606170654
8'b00001101,  // 0.8414360880851746
8'b00000110,  // 0.397830605506897
8'b00000110,  // 0.4105983078479767
8'b11000101,  // -3.657735586166382
8'b11110001,  // -0.8977976441383362
8'b00011011,  // 1.7051936388015747
8'b11101011,  // -1.2765135765075684
8'b11110110,  // -0.5837795734405518
8'b00101011,  // 2.699671983718872
8'b00000011,  // 0.2170683741569519
8'b00001110,  // 0.8814588785171509
8'b11010101,  // -2.634300947189331
8'b11100001,  // -1.877297282218933
8'b00011010,  // 1.6625694036483765
8'b00101011,  // 2.7459704875946045
8'b11111000,  // -0.47838035225868225
8'b00011011,  // 1.6984987258911133
8'b00001101,  // 0.8548859357833862
8'b00010000,  // 1.0045719146728516
8'b00010110,  // 1.4197649955749512
8'b00001101,  // 0.832463800907135
8'b00001000,  // 0.5434179306030273
8'b00001110,  // 0.9277304410934448
8'b11111010,  // -0.3426123857498169
8'b11110111,  // -0.5587119460105896
8'b11110110,  // -0.6208624839782715
8'b11101011,  // -1.2802538871765137
8'b00000000,  // 0.05940237268805504
8'b11110010,  // -0.8213341236114502
8'b00001110,  // 0.8783953189849854
8'b11110000   // -0.949700653553009
};
endpackage