// Width: 16
// NFRAC: 6
package dense_1_16_6;

localparam logic signed [15:0] weights [16][64] = '{ 
{16'b0000000000010000, 16'b1111111111010110, 16'b1111111111110100, 16'b1111111111110001, 16'b1111111111100110, 16'b0000000000000111, 16'b1111111110111101, 16'b0000000000000000, 16'b0000000000000011, 16'b0000000000010000, 16'b0000000000000000, 16'b1111111111100110, 16'b1111111111111111, 16'b0000000000001101, 16'b0000000000000010, 16'b1111111111101111, 16'b0000000000001110, 16'b0000000000000011, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000011000, 16'b1111111111101010, 16'b1111111111111110, 16'b0000000000011110, 16'b1111111111101011, 16'b1111111111010100, 16'b1111111111101110, 16'b1111111111110011, 16'b1111111111111001, 16'b1111111111111111, 16'b0000000000000010, 16'b0000000000001111, 16'b0000000000001100, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000010011, 16'b1111111111111110, 16'b1111111111101111, 16'b0000000000000001, 16'b0000000000001100, 16'b1111111111111111, 16'b0000000000010001, 16'b1111111111101110, 16'b0000000000111011, 16'b1111111111111111, 16'b0000000000011100, 16'b0000000000000000, 16'b0000000000001011, 16'b0000000000001100, 16'b1111111111111110, 16'b0000000000000000, 16'b0000000000001010, 16'b0000000000001101, 16'b0000000000000100, 16'b1111111111111000, 16'b1111111111101100, 16'b0000000000100010, 16'b1111111111100000, 16'b0000000000011101, 16'b1111111111101001, 16'b0000000000110010, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000101}, 
{16'b0000000000000000, 16'b1111111111101011, 16'b1111111111110111, 16'b1111111111101110, 16'b1111111111101011, 16'b0000000000000110, 16'b1111111111001111, 16'b1111111111111111, 16'b1111111111110001, 16'b0000000000001011, 16'b0000000000000000, 16'b1111111111111010, 16'b0000000000001100, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000001101, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111110100, 16'b1111111111101111, 16'b0000000000011100, 16'b1111111111111010, 16'b0000000000000011, 16'b0000000000101100, 16'b0000000000010000, 16'b1111111111110001, 16'b1111111111110001, 16'b1111111111111111, 16'b1111111111111001, 16'b1111111111100110, 16'b1111111111111100, 16'b0000000000011101, 16'b0000000000010001, 16'b0000000000100011, 16'b0000000000101000, 16'b0000000000000011, 16'b1111111111111000, 16'b1111111111100100, 16'b0000000000000011, 16'b0000000000001100, 16'b0000000000000001, 16'b0000000000001101, 16'b1111111111110010, 16'b0000000000010000, 16'b0000000000001011, 16'b0000000000000011, 16'b1111111111101010, 16'b0000000000000101, 16'b0000000000010000, 16'b0000000000000001, 16'b0000000000000001, 16'b0000000001001010, 16'b1111111111111011, 16'b1111111111111001, 16'b1111111111111100, 16'b1111111111111111, 16'b0000000000010000, 16'b1111111111101000, 16'b0000000000111111, 16'b0000000000000000, 16'b0000000000100001, 16'b0000000000001111, 16'b0000000000110100, 16'b0000000000001001}, 
{16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111010, 16'b1111111111110100, 16'b1111111111110100, 16'b0000000000000010, 16'b0000000001011110, 16'b1111111111111111, 16'b1111111110101110, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111110, 16'b1111111111110001, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000001010, 16'b0000000000111001, 16'b1111111111111111, 16'b0000000000000100, 16'b0000000000000000, 16'b0000000000011010, 16'b1111111111010001, 16'b0000000000100100, 16'b1111111111010010, 16'b0000000000111100, 16'b1111111111101001, 16'b1111111111110000, 16'b1111111111010010, 16'b0000000001010001, 16'b0000000000010001, 16'b0000000000000000, 16'b0000000000100001, 16'b0000000001000001, 16'b1111111110110011, 16'b1111111111111001, 16'b0000000000000010, 16'b1111111111110001, 16'b0000000000111001, 16'b1111111111111101, 16'b0000000000010100, 16'b0000000000010101, 16'b0000000000010111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111110, 16'b0000000000001010, 16'b1111111111101110, 16'b1111111111110101, 16'b1111111111111110, 16'b0000000000011001, 16'b1111111111110100, 16'b0000000000001001, 16'b1111111111111111, 16'b0000000000001000, 16'b1111111111110100, 16'b1111111111111111, 16'b1111111111101100, 16'b1111111111010101, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000001100010, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111101100}, 
{16'b1111111111100010, 16'b1111111111101000, 16'b1111111111010011, 16'b0000000000010011, 16'b1111111111101011, 16'b1111111110101001, 16'b1111111111111000, 16'b1111111111101100, 16'b0000000000001110, 16'b1111111111111111, 16'b0000000001010000, 16'b1111111111111001, 16'b1111111111001101, 16'b0000000000100101, 16'b0000000000000001, 16'b1111111111111111, 16'b1111111111100011, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111110001, 16'b1111111110110110, 16'b1111111111111000, 16'b1111111111010011, 16'b0000000000001100, 16'b1111111111100111, 16'b1111111111000101, 16'b0000000000010100, 16'b0000000000101111, 16'b0000000001010010, 16'b1111111111100010, 16'b1111111111011010, 16'b0000000000000100, 16'b0000000000100000, 16'b1111111111001010, 16'b1111111111101011, 16'b0000000000000000, 16'b1111111111010001, 16'b0000000000001111, 16'b1111111111100011, 16'b0000000000000111, 16'b0000000000011101, 16'b0000000000001010, 16'b0000000000000000, 16'b0000000000000001, 16'b0000000000100011, 16'b1111111111110011, 16'b1111111111111111, 16'b1111111111101001, 16'b1111111111111111, 16'b1111111111111001, 16'b1111111111011000, 16'b0000000000000101, 16'b1111111111111111, 16'b0000000000001101, 16'b0000000000010100, 16'b0000000000101001, 16'b1111111111000010, 16'b1111111111000100, 16'b1111111111010010, 16'b0000000000110111, 16'b0000000001101111, 16'b1111111111000110, 16'b1111111111111100, 16'b0000000000011011}, 
{16'b0000000000010101, 16'b1111111111011000, 16'b1111111111101111, 16'b1111111111111111, 16'b1111111111110110, 16'b0000000000010101, 16'b0000000000001100, 16'b1111111111111111, 16'b1111111111011001, 16'b1111111111110000, 16'b1111111111101000, 16'b0000000000000011, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111101, 16'b0000000000010110, 16'b0000000000001000, 16'b1111111111100110, 16'b0000000000000001, 16'b0000000000000000, 16'b0000000000001101, 16'b1111111111111000, 16'b0000000000000100, 16'b1111111111111110, 16'b0000000001000100, 16'b1111111111110100, 16'b1111111111101110, 16'b1111111111100110, 16'b0000000000000000, 16'b0000000000001010, 16'b0000000000000111, 16'b0000000000010001, 16'b1111111111111111, 16'b0000000000000100, 16'b0000000000001000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000111000, 16'b1111111111101101, 16'b1111111111111011, 16'b0000000000011011, 16'b0000000000001111, 16'b1111111111100000, 16'b0000000000000000, 16'b1111111110111011, 16'b1111111111111111, 16'b1111111111111000, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111110, 16'b1111111111111111, 16'b0000000000001100, 16'b1111111111111111, 16'b0000000000010100, 16'b1111111111110011, 16'b1111111111010000, 16'b1111111111100010, 16'b1111111111011111, 16'b1111111111011000, 16'b0000000000101111, 16'b0000000001010111, 16'b0000000000110010, 16'b0000000000000111, 16'b1111111111111111}, 
{16'b1111111111100011, 16'b1111111111010111, 16'b0000000000000000, 16'b0000000000010011, 16'b0000000000010010, 16'b1111111111110010, 16'b0000000000100101, 16'b1111111111111111, 16'b0000000000001111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111011, 16'b1111111111110100, 16'b0000000000100101, 16'b1111111111111010, 16'b0000000000000000, 16'b1111111111011000, 16'b1111111111101001, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111100, 16'b1111111111101011, 16'b1111111111101011, 16'b0000000000011101, 16'b1111111111101011, 16'b1111111111111111, 16'b0000000000010000, 16'b1111111111111011, 16'b1111111111000100, 16'b1111111111111111, 16'b1111111111111011, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000010, 16'b0000000000001000, 16'b0000000000010110, 16'b0000000000000000, 16'b1111111111111001, 16'b1111111111101111, 16'b1111111111111111, 16'b1111111111110101, 16'b1111111111011110, 16'b0000000000011001, 16'b0000000000000000, 16'b0000000000100110, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000110, 16'b1111111111100101, 16'b0000000000001110, 16'b0000000000000000, 16'b1111111111111001, 16'b1111111111101000, 16'b0000000000011000, 16'b1111111111111111, 16'b0000000000010110, 16'b0000000000001101, 16'b0000000000001101, 16'b1111111111111110, 16'b1111111111111111, 16'b1111111111001100, 16'b1111111111110111, 16'b1111111111111100, 16'b1111111111111111}, 
{16'b1111111111101101, 16'b1111111111101010, 16'b1111111111100100, 16'b1111111111111011, 16'b1111111111110111, 16'b0000000000000110, 16'b1111111111010011, 16'b1111111111110110, 16'b1111111111110001, 16'b1111111111111111, 16'b1111111111101101, 16'b0000000000010110, 16'b0000000000000010, 16'b0000000000001000, 16'b0000000000010011, 16'b0000000000000000, 16'b0000000000110011, 16'b0000000000000101, 16'b0000000000001111, 16'b0000000000010001, 16'b1111111111110101, 16'b0000000000010111, 16'b1111111111110000, 16'b1111111111011111, 16'b0000000000001011, 16'b0000000000100001, 16'b1111111111111111, 16'b0000000000000011, 16'b1111111111000011, 16'b0000000000010010, 16'b0000000000010001, 16'b1111111111101000, 16'b0000000000011110, 16'b0000000000101010, 16'b0000000000000000, 16'b0000000000010101, 16'b1111111111111111, 16'b0000000000010010, 16'b0000000000001100, 16'b0000000000000000, 16'b1111111111111000, 16'b1111111111101000, 16'b0000000000001001, 16'b0000000000011110, 16'b0000000000100001, 16'b1111111111110101, 16'b1111111111111010, 16'b1111111111110011, 16'b1111111111110111, 16'b0000000000000111, 16'b0000000000000000, 16'b0000000000000010, 16'b0000000000000000, 16'b0000000000001011, 16'b1111111111110100, 16'b0000000000110001, 16'b0000000000010110, 16'b1111111111111110, 16'b0000000000011000, 16'b0000000000001101, 16'b1111111110010111, 16'b1111111111011011, 16'b1111111111110100, 16'b1111111111111111}, 
{16'b0000000000000000, 16'b0000000000001111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111101011, 16'b1111111111111110, 16'b1111111111101111, 16'b0000000000000000, 16'b0000000000000001, 16'b0000000000011000, 16'b0000000000000000, 16'b1111111111100111, 16'b1111111111111011, 16'b0000000000000000, 16'b1111111111111100, 16'b1111111111100011, 16'b1111111111001001, 16'b1111111111111111, 16'b1111111111011001, 16'b1111111111100011, 16'b1111111111100111, 16'b0000000000010110, 16'b0000000000000011, 16'b1111111111110110, 16'b1111111111100100, 16'b0000000000001001, 16'b0000000000000000, 16'b0000000000011111, 16'b0000000000110011, 16'b1111111111111101, 16'b0000000000000000, 16'b0000000000001110, 16'b1111111111010100, 16'b1111111111101000, 16'b0000000000000011, 16'b0000000000000101, 16'b1111111111101110, 16'b0000000000001111, 16'b0000000000001000, 16'b1111111111110110, 16'b1111111111100101, 16'b1111111111111101, 16'b0000000000000010, 16'b1111111111110101, 16'b0000000000000011, 16'b0000000000001110, 16'b1111111111111000, 16'b0000000000000001, 16'b0000000000000000, 16'b1111111111110010, 16'b1111111111100111, 16'b0000000000011010, 16'b0000000000001000, 16'b1111111111110100, 16'b0000000000001000, 16'b1111111111111100, 16'b1111111111100001, 16'b1111111111110111, 16'b1111111111111100, 16'b1111111111111011, 16'b0000000000110101, 16'b0000000000001100, 16'b1111111111111100, 16'b1111111111111111}, 
{16'b0000000000000000, 16'b0000000000100101, 16'b1111111111011010, 16'b1111111111110001, 16'b0000000000010100, 16'b1111111111110010, 16'b0000000001001101, 16'b1111111111101101, 16'b1111111111111111, 16'b0000000000010010, 16'b0000000000010000, 16'b1111111111111111, 16'b1111111111111100, 16'b1111111111100001, 16'b0000000000010010, 16'b0000000000001010, 16'b1111111111110011, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000010000, 16'b1111111111100010, 16'b0000000000011001, 16'b0000000000100111, 16'b1111111111111010, 16'b1111111111111111, 16'b1111111111111110, 16'b1111111111111111, 16'b0000000000101111, 16'b0000000000000000, 16'b1111111111101110, 16'b0000000000000000, 16'b0000000000011000, 16'b1111111111001100, 16'b1111111111011101, 16'b0000000000001100, 16'b0000000000001000, 16'b1111111111011011, 16'b1111111111110011, 16'b1111111111110010, 16'b0000000000011001, 16'b0000000000011001, 16'b0000000000000000, 16'b1111111111101110, 16'b0000000000000000, 16'b0000000000011001, 16'b1111111111111100, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000001111, 16'b1111111111111100, 16'b1111111111110011, 16'b0000000000010110, 16'b1111111111110010, 16'b0000000000010001, 16'b0000000000100101, 16'b0000000000000010, 16'b0000000000010000, 16'b1111111111100110, 16'b1111111111101000, 16'b0000000000110101, 16'b1111111111110111, 16'b0000000000000010, 16'b1111111111111010}, 
{16'b0000000000000001, 16'b1111111111100011, 16'b0000000000010111, 16'b1111111111101101, 16'b1111111111111111, 16'b0000000000001101, 16'b1111111111011010, 16'b0000000000001100, 16'b0000000000011111, 16'b0000000000001001, 16'b0000000000010111, 16'b0000000000010100, 16'b1111111111101100, 16'b1111111111111011, 16'b1111111111111100, 16'b0000000000000000, 16'b1111111111000010, 16'b0000000000010100, 16'b1111111111111101, 16'b0000000000000001, 16'b1111111111101001, 16'b0000000000000100, 16'b0000000000001001, 16'b1111111111111111, 16'b1111111111100010, 16'b1111111111111100, 16'b1111111111111010, 16'b0000000001001111, 16'b1111111111010101, 16'b0000000000000100, 16'b0000000000000110, 16'b1111111111111100, 16'b1111111111110001, 16'b0000000000000111, 16'b1111111111111010, 16'b1111111111110111, 16'b1111111111110100, 16'b1111111111110010, 16'b1111111111111110, 16'b1111111111101100, 16'b0000000000010100, 16'b0000000000000111, 16'b0000000000011111, 16'b0000000000000101, 16'b0000000000000010, 16'b1111111111101101, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000001100, 16'b0000000000001011, 16'b0000000000010010, 16'b1111111111111111, 16'b1111111111101101, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000010100, 16'b1111111111110011, 16'b1111111111011100, 16'b0000000000100011, 16'b1111111111101101, 16'b0000000001001010, 16'b1111111111111110, 16'b1111111111101001}, 
{16'b1111111111011011, 16'b1111111111111111, 16'b1111111111100101, 16'b0000000000001110, 16'b0000000000010000, 16'b1111111111111001, 16'b0000000000100001, 16'b1111111111110101, 16'b1111111111100001, 16'b1111111111101000, 16'b1111111111101111, 16'b1111111111100001, 16'b1111111111110001, 16'b0000000000001100, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000110101, 16'b1111111111111101, 16'b1111111111111111, 16'b0000000000011010, 16'b0000000000010010, 16'b1111111111011010, 16'b1111111111100111, 16'b0000000000001100, 16'b1111111111100100, 16'b1111111111111110, 16'b1111111111101111, 16'b1111111111101010, 16'b1111111111100100, 16'b0000000000010011, 16'b0000000000001110, 16'b1111111111110110, 16'b1111111111111011, 16'b1111111111000001, 16'b1111111111110100, 16'b0000000000000011, 16'b1111111111110111, 16'b1111111111101101, 16'b1111111111111111, 16'b0000000000000111, 16'b1111111111111000, 16'b1111111111111111, 16'b1111111111111101, 16'b1111111111010101, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000010101, 16'b1111111111111000, 16'b0000000000011011, 16'b1111111111110011, 16'b0000000000010010, 16'b1111111111111111, 16'b0000000000001110, 16'b1111111111100110, 16'b1111111111111111, 16'b0000000000100000, 16'b0000000000010100, 16'b0000000000010010, 16'b0000000000000001, 16'b1111111111100110, 16'b1111111111101100, 16'b1111111111010100, 16'b1111111111111111, 16'b0000000000000110}, 
{16'b0000000000010011, 16'b0000000000000000, 16'b0000000000001000, 16'b1111111111111111, 16'b0000000000001001, 16'b1111111111110111, 16'b0000000000001111, 16'b0000000000000010, 16'b0000000000001000, 16'b0000000000010101, 16'b1111111111101111, 16'b1111111111111110, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111010101, 16'b1111111111101100, 16'b0000000000101000, 16'b1111111111111110, 16'b1111111111111100, 16'b0000000000000000, 16'b1111111111100111, 16'b0000000000000000, 16'b0000000000010000, 16'b0000000000000010, 16'b0000000000000010, 16'b0000000000010101, 16'b0000000000000000, 16'b0000000000000010, 16'b0000000000000000, 16'b1111111111111100, 16'b1111111111110011, 16'b1111111111010101, 16'b0000000000010000, 16'b0000000000010101, 16'b1111111111111110, 16'b1111111111110000, 16'b0000000000000000, 16'b1111111111010110, 16'b1111111111111101, 16'b1111111111111111, 16'b0000000000001100, 16'b1111111111110111, 16'b1111111111111111, 16'b0000000000110110, 16'b0000000000011100, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111110000, 16'b0000000000001001, 16'b0000000000001001, 16'b0000000000001011, 16'b0000000000001010, 16'b0000000000011000, 16'b0000000000010110, 16'b0000000000101010, 16'b1111111111110111, 16'b0000000000011001, 16'b0000000000001001, 16'b1111111111101011, 16'b0000000000000111, 16'b1111111111100111, 16'b1111111111100011, 16'b1111111111100000}, 
{16'b0000000000000000, 16'b0000000000001110, 16'b1111111111110011, 16'b0000000000000000, 16'b1111111111111100, 16'b1111111111111101, 16'b1111111111010101, 16'b1111111111111111, 16'b0000000000010000, 16'b0000000000001111, 16'b0000000000001111, 16'b1111111111100110, 16'b1111111111111010, 16'b0000000000010010, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111001010, 16'b1111111111111111, 16'b0000000000010111, 16'b0000000000000100, 16'b0000000000001111, 16'b1111111111111000, 16'b0000000000001111, 16'b0000000000011001, 16'b1111111111101001, 16'b1111111111101110, 16'b1111111111111111, 16'b1111111111111010, 16'b0000000000000100, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000010100, 16'b1111111111010000, 16'b0000000000010111, 16'b0000000000100000, 16'b0000000000000111, 16'b0000000000000111, 16'b1111111111111001, 16'b0000000000000111, 16'b1111111111111001, 16'b1111111111101111, 16'b1111111111111100, 16'b0000000000001010, 16'b0000000000101100, 16'b1111111111001001, 16'b1111111111100011, 16'b0000000000001100, 16'b1111111111111001, 16'b0000000000011100, 16'b1111111111110000, 16'b1111111111101010, 16'b1111111111101110, 16'b1111111111111111, 16'b0000000000000111, 16'b1111111111110101, 16'b1111111111001010, 16'b1111111111110110, 16'b1111111111111111, 16'b0000000000000010, 16'b1111111111011000, 16'b0000000001000111, 16'b1111111111011101, 16'b0000000000100010, 16'b0000000000001001}, 
{16'b0000000000000101, 16'b1111111111110011, 16'b0000000000101000, 16'b1111111111101100, 16'b1111111111100010, 16'b0000000000000101, 16'b0000000000010011, 16'b0000000000010011, 16'b1111111111110100, 16'b1111111111110101, 16'b0000000000000011, 16'b0000000000001110, 16'b0000000000001111, 16'b0000000000000011, 16'b1111111111110010, 16'b0000000000001000, 16'b0000000000011110, 16'b1111111111111111, 16'b1111111111101110, 16'b0000000000000000, 16'b0000000000000100, 16'b0000000000000001, 16'b1111111111101101, 16'b0000000000000111, 16'b0000000000110010, 16'b0000000000000000, 16'b0000000000001011, 16'b1111111111001101, 16'b1111111111111011, 16'b0000000000000000, 16'b1111111111110011, 16'b1111111111101100, 16'b0000000000011101, 16'b1111111111111110, 16'b1111111111111101, 16'b1111111111101100, 16'b0000000000001000, 16'b0000000000010010, 16'b1111111111111111, 16'b1111111111111101, 16'b1111111111110100, 16'b0000000000001110, 16'b0000000000000000, 16'b1111111111010100, 16'b0000000000010011, 16'b0000000000011001, 16'b1111111111111111, 16'b0000000000000001, 16'b1111111111100100, 16'b1111111111111011, 16'b1111111111111111, 16'b1111111111101011, 16'b0000000000000000, 16'b1111111111110100, 16'b0000000000000011, 16'b1111111111001011, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000010001, 16'b0000000000100100, 16'b1111111111010011, 16'b0000000000100001, 16'b0000000000000010, 16'b1111111111111011}, 
{16'b0000000000010010, 16'b0000000001001111, 16'b0000000000011111, 16'b0000000000010010, 16'b1111111111100001, 16'b1111111111101011, 16'b1111111101011001, 16'b1111111111100010, 16'b0000000000011001, 16'b1111111111111111, 16'b0000000000010010, 16'b0000000000110111, 16'b0000000000000100, 16'b0000000000000000, 16'b1111111111111110, 16'b0000000000000000, 16'b1111111111110011, 16'b1111111111110011, 16'b0000000000001110, 16'b1111111111011111, 16'b1111111111010101, 16'b1111111111111001, 16'b1111111111011010, 16'b0000000000000001, 16'b1111111101101110, 16'b0000000000110100, 16'b0000000000111111, 16'b0000000000100110, 16'b1111111110010000, 16'b1111111111101011, 16'b1111111111010011, 16'b1111111111001010, 16'b1111111101011110, 16'b0000000000101011, 16'b1111111111111101, 16'b0000000000010100, 16'b0000000000000001, 16'b1111111110100100, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000010, 16'b0000000001000001, 16'b1111111111110010, 16'b1111111111010110, 16'b0000000000111001, 16'b1111111111100011, 16'b1111111111101011, 16'b1111111111100110, 16'b0000000000011110, 16'b0000000000100010, 16'b1111111111111011, 16'b1111111111101001, 16'b1111111111111111, 16'b1111111111111000, 16'b0000000000000000, 16'b1111111111100111, 16'b0000000000100110, 16'b0000000001000101, 16'b0000000000101101, 16'b1111111111000101, 16'b1111111100010011, 16'b0000000000111000, 16'b0000000000000101, 16'b0000000000010100}, 
{16'b1111111111110000, 16'b0000000000010101, 16'b0000000000010100, 16'b1111111111111111, 16'b1111111111101000, 16'b1111111111111010, 16'b1111111111100111, 16'b1111111111111100, 16'b0000000000001001, 16'b1111111111111011, 16'b1111111111111110, 16'b1111111111111101, 16'b1111111111111111, 16'b1111111111110100, 16'b1111111111111110, 16'b1111111111111001, 16'b0000000000010100, 16'b1111111111111111, 16'b1111111111010110, 16'b0000000000011101, 16'b0000000000100110, 16'b0000000000011010, 16'b1111111111101011, 16'b1111111111110111, 16'b1111111111101001, 16'b1111111111101101, 16'b0000000000001110, 16'b0000000000001110, 16'b0000000000001110, 16'b0000000000010111, 16'b0000000000000010, 16'b0000000000011000, 16'b1111111111111101, 16'b0000000000000000, 16'b0000000000010011, 16'b0000000000001000, 16'b1111111111111011, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111101101, 16'b1111111111110001, 16'b1111111111111000, 16'b1111111111101001, 16'b0000000000011100, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111010, 16'b1111111111110110, 16'b1111111111001100, 16'b1111111111111101, 16'b1111111111110001, 16'b1111111111110110, 16'b1111111111111001, 16'b0000000000010000, 16'b0000000000101011, 16'b0000000000001011, 16'b1111111111111111, 16'b1111111111101010, 16'b1111111111111110, 16'b0000000000000000, 16'b0000000000010100, 16'b1111111111111110, 16'b0000000000000010, 16'b0000000000000000}
};

localparam logic signed [15:0] bias [64] = '{
16'b1111111111111101,  // -0.037350185215473175
16'b0000000000010001,  // 0.27355897426605225
16'b1111111111111000,  // -0.12378914654254913
16'b1111111111111011,  // -0.064457006752491
16'b0000000000000011,  // 0.05452875792980194
16'b0000000000000111,  // 0.11671770364046097
16'b0000000000001000,  // 0.13640816509723663
16'b0000000000000100,  // 0.07482525706291199
16'b0000000000000010,  // 0.04674031585454941
16'b1111111111110011,  // -0.20146161317825317
16'b1111111111111001,  // -0.09910125285387039
16'b0000000000001001,  // 0.15104414522647858
16'b1111111111111001,  // -0.10221704095602036
16'b1111111111110110,  // -0.1461549550294876
16'b1111111111111010,  // -0.08641516417264938
16'b0000000000001010,  // 0.16613510251045227
16'b1111111111111010,  // -0.0836295336484909
16'b1111111111111100,  // -0.05756539851427078
16'b1111111111111101,  // -0.03229188174009323
16'b1111111111111110,  // -0.028388574719429016
16'b0000000000001000,  // 0.1260243058204651
16'b1111111111111101,  // -0.037064336240291595
16'b0000000000001100,  // 0.19336333870887756
16'b0000000000000001,  // 0.02124214917421341
16'b0000000000011111,  // 0.4985624849796295
16'b0000000000000001,  // 0.0158411655575037
16'b1111111111111010,  // -0.08296407759189606
16'b0000000000000111,  // 0.11056788265705109
16'b0000000000000000,  // 0.01173810102045536
16'b1111111111111001,  // -0.10843746364116669
16'b0000000000010001,  // 0.27439257502555847
16'b0000000000000101,  // 0.09199801832437515
16'b0000000000010001,  // 0.27419957518577576
16'b0000000000010001,  // 0.27063727378845215
16'b1111111111110000,  // -0.24828937649726868
16'b0000000000000101,  // 0.07818280160427094
16'b1111111111111111,  // -0.005749030504375696
16'b0000000000000110,  // 0.10850494354963303
16'b0000000000001000,  // 0.13591453433036804
16'b1111111111111000,  // -0.12088628858327866
16'b1111111111111100,  // -0.05666546896100044
16'b0000000000000101,  // 0.09311636537313461
16'b0000000000000011,  // 0.05477767437696457
16'b0000000000000001,  // 0.029585206881165504
16'b1111111111101100,  // -0.31209176778793335
16'b1111111111111010,  // -0.08465463668107986
16'b1111111111110101,  // -0.16775836050510406
16'b0000000000001001,  // 0.14762157201766968
16'b1111111111110000,  // -0.23618532717227936
16'b0000000000000100,  // 0.06535740196704865
16'b1111111111110111,  // -0.12853026390075684
16'b1111111111110111,  // -0.13802281022071838
16'b1111111111110110,  // -0.15156887471675873
16'b0000000000000101,  // 0.07979883998632431
16'b0000000000001011,  // 0.18141601979732513
16'b1111111111111100,  // -0.054039113223552704
16'b1111111111111111,  // -0.010052933357656002
16'b0000000000000100,  // 0.06611225008964539
16'b0000000000000011,  // 0.05053366720676422
16'b0000000000000001,  // 0.026860840618610382
16'b0000000000000010,  // 0.03283466026186943
16'b0000000000001001,  // 0.15558314323425293
16'b1111111111101101,  // -0.2863388657569885
16'b1111111111111010   // -0.08769102394580841
};
endpackage