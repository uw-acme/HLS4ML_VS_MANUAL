// Width: 13
// NFRAC: 6
package dense_4_13_6;

localparam logic signed [12:0] weights [32][5] = '{ 
{13'b1111111111111, 13'b0000000010100, 13'b1111111101100, 13'b0000000000100, 13'b1111111111001}, 
{13'b1111111011100, 13'b1111111111100, 13'b0000000011101, 13'b1111111111111, 13'b0000000000001}, 
{13'b0000000010111, 13'b0000000001101, 13'b1111111111110, 13'b1111111100110, 13'b1111111110010}, 
{13'b1111111100111, 13'b1111111101000, 13'b1111111111000, 13'b0000000010011, 13'b0000000001111}, 
{13'b0000000000111, 13'b0000000001000, 13'b0000000001010, 13'b1111111111110, 13'b1111110111111}, 
{13'b0000000010100, 13'b1111111100110, 13'b0000000001011, 13'b1111111110101, 13'b1111111110101}, 
{13'b1111111100110, 13'b0000000000010, 13'b1111111111111, 13'b0000000001011, 13'b0000000000100}, 
{13'b1111111111111, 13'b0000000010010, 13'b1111111100110, 13'b0000000001010, 13'b0000000001000}, 
{13'b0000000001010, 13'b1111111110101, 13'b0000000000000, 13'b1111111100010, 13'b1111111110000}, 
{13'b1111111111111, 13'b1111111101110, 13'b0000000001011, 13'b0000000011011, 13'b0000000000000}, 
{13'b1111111110111, 13'b1111111110110, 13'b0000000000000, 13'b0000000100101, 13'b1111111101110}, 
{13'b0000000001010, 13'b0000000001110, 13'b1111111101010, 13'b1111111111110, 13'b0000000000111}, 
{13'b0000000000000, 13'b0000000001010, 13'b0000000000000, 13'b1111111110010, 13'b1111111011000}, 
{13'b0000000001011, 13'b0000000000100, 13'b0000000011010, 13'b1111111111011, 13'b1111111100100}, 
{13'b0000000000101, 13'b1111111111100, 13'b1111111101000, 13'b1111111111101, 13'b0000000100010}, 
{13'b1111111100001, 13'b1111111110000, 13'b1111111110001, 13'b0000000011001, 13'b0000000000010}, 
{13'b0000000010110, 13'b1111111110101, 13'b1111111110111, 13'b1111111110001, 13'b1111111111100}, 
{13'b0000000001100, 13'b1111111111101, 13'b1111111100101, 13'b1111111111110, 13'b0000000000100}, 
{13'b0000000010000, 13'b0000000000010, 13'b1111111110010, 13'b0000000000000, 13'b1111111100111}, 
{13'b0000000001110, 13'b1111111111010, 13'b1111111110010, 13'b0000000001101, 13'b0000000000110}, 
{13'b0000000000100, 13'b1111111111110, 13'b0000000010011, 13'b1111111100100, 13'b1111111111110}, 
{13'b0000000000000, 13'b0000000000111, 13'b0000000011111, 13'b1111111011110, 13'b1111111011000}, 
{13'b1111111111001, 13'b0000000000111, 13'b0000000001011, 13'b1111111101001, 13'b0000000100001}, 
{13'b1111111111111, 13'b0000000001010, 13'b0000000010010, 13'b0000000000010, 13'b1111111011011}, 
{13'b1111111110101, 13'b0000000010111, 13'b1111111110001, 13'b0000000000000, 13'b0000000011000}, 
{13'b0000000000001, 13'b0000000010001, 13'b0000000000001, 13'b1111111010000, 13'b0000000100011}, 
{13'b1111111100010, 13'b1111111110000, 13'b0000000001101, 13'b0000000001111, 13'b0000000001100}, 
{13'b0000000000000, 13'b0000000001111, 13'b1111111111101, 13'b1111111110110, 13'b0000000000010}, 
{13'b1111111111001, 13'b0000000001111, 13'b1111111011111, 13'b0000000001000, 13'b1111111110101}, 
{13'b1111111111110, 13'b0000000001001, 13'b1111111110101, 13'b1111111100110, 13'b0000000100101}, 
{13'b0000000011100, 13'b0000000000100, 13'b0000000010100, 13'b1111111011010, 13'b1111111101011}, 
{13'b1111111111100, 13'b1111111100111, 13'b0000000010111, 13'b0000000000100, 13'b0000000001000}
};

localparam logic signed [12:0] bias [5] = '{
13'b1111111111100,  // -0.06223141402006149
13'b1111111111011,  // -0.06270556896924973
13'b1111111111011,  // -0.07014333456754684
13'b0000000000101,  // 0.0820775106549263
13'b0000000001101   // 0.2155742198228836
};
endpackage