// Width: 10
// NFRAC: 5
package dense_4_10_5;

localparam logic signed [9:0] weights [32][5] = '{ 
{10'b1111111111, 10'b0000001010, 10'b1111110110, 10'b0000000010, 10'b1111111100}, 
{10'b1111101110, 10'b1111111110, 10'b0000001110, 10'b1111111111, 10'b0000000000}, 
{10'b0000001011, 10'b0000000110, 10'b1111111111, 10'b1111110011, 10'b1111111001}, 
{10'b1111110011, 10'b1111110100, 10'b1111111100, 10'b0000001001, 10'b0000000111}, 
{10'b0000000011, 10'b0000000100, 10'b0000000101, 10'b1111111111, 10'b1111011111}, 
{10'b0000001010, 10'b1111110011, 10'b0000000101, 10'b1111111010, 10'b1111111010}, 
{10'b1111110011, 10'b0000000001, 10'b1111111111, 10'b0000000101, 10'b0000000010}, 
{10'b1111111111, 10'b0000001001, 10'b1111110011, 10'b0000000101, 10'b0000000100}, 
{10'b0000000101, 10'b1111111010, 10'b0000000000, 10'b1111110001, 10'b1111111000}, 
{10'b1111111111, 10'b1111110111, 10'b0000000101, 10'b0000001101, 10'b0000000000}, 
{10'b1111111011, 10'b1111111011, 10'b0000000000, 10'b0000010010, 10'b1111110111}, 
{10'b0000000101, 10'b0000000111, 10'b1111110101, 10'b1111111111, 10'b0000000011}, 
{10'b0000000000, 10'b0000000101, 10'b0000000000, 10'b1111111001, 10'b1111101100}, 
{10'b0000000101, 10'b0000000010, 10'b0000001101, 10'b1111111101, 10'b1111110010}, 
{10'b0000000010, 10'b1111111110, 10'b1111110100, 10'b1111111110, 10'b0000010001}, 
{10'b1111110000, 10'b1111111000, 10'b1111111000, 10'b0000001100, 10'b0000000001}, 
{10'b0000001011, 10'b1111111010, 10'b1111111011, 10'b1111111000, 10'b1111111110}, 
{10'b0000000110, 10'b1111111110, 10'b1111110010, 10'b1111111111, 10'b0000000010}, 
{10'b0000001000, 10'b0000000001, 10'b1111111001, 10'b0000000000, 10'b1111110011}, 
{10'b0000000111, 10'b1111111101, 10'b1111111001, 10'b0000000110, 10'b0000000011}, 
{10'b0000000010, 10'b1111111111, 10'b0000001001, 10'b1111110010, 10'b1111111111}, 
{10'b0000000000, 10'b0000000011, 10'b0000001111, 10'b1111101111, 10'b1111101100}, 
{10'b1111111100, 10'b0000000011, 10'b0000000101, 10'b1111110100, 10'b0000010000}, 
{10'b1111111111, 10'b0000000101, 10'b0000001001, 10'b0000000001, 10'b1111101101}, 
{10'b1111111010, 10'b0000001011, 10'b1111111000, 10'b0000000000, 10'b0000001100}, 
{10'b0000000000, 10'b0000001000, 10'b0000000000, 10'b1111101000, 10'b0000010001}, 
{10'b1111110001, 10'b1111111000, 10'b0000000110, 10'b0000000111, 10'b0000000110}, 
{10'b0000000000, 10'b0000000111, 10'b1111111110, 10'b1111111011, 10'b0000000001}, 
{10'b1111111100, 10'b0000000111, 10'b1111101111, 10'b0000000100, 10'b1111111010}, 
{10'b1111111111, 10'b0000000100, 10'b1111111010, 10'b1111110011, 10'b0000010010}, 
{10'b0000001110, 10'b0000000010, 10'b0000001010, 10'b1111101101, 10'b1111110101}, 
{10'b1111111110, 10'b1111110011, 10'b0000001011, 10'b0000000010, 10'b0000000100}
};

localparam logic signed [9:0] bias [5] = '{
10'b1111111110,  // -0.06223141402006149
10'b1111111101,  // -0.06270556896924973
10'b1111111101,  // -0.07014333456754684
10'b0000000010,  // 0.0820775106549263
10'b0000000110   // 0.2155742198228836
};
endpackage