// Width: 17
// NFRAC: 8
package dense_4_17_8;

localparam logic signed [16:0] weights [32][5] = '{ 
{17'b11111111111111100, 17'b00000000001010000, 17'b11111111110110011, 17'b00000000000010000, 17'b11111111111100100}, 
{17'b11111111101110001, 17'b11111111111110001, 17'b00000000001110101, 17'b11111111111111100, 17'b00000000000000100}, 
{17'b00000000001011111, 17'b00000000000110110, 17'b11111111111111000, 17'b11111111110011000, 17'b11111111111001010}, 
{17'b11111111110011111, 17'b11111111110100000, 17'b11111111111100011, 17'b00000000001001110, 17'b00000000000111100}, 
{17'b00000000000011111, 17'b00000000000100000, 17'b00000000000101000, 17'b11111111111111011, 17'b11111111011111100}, 
{17'b00000000001010011, 17'b11111111110011011, 17'b00000000000101110, 17'b11111111111010110, 17'b11111111111010100}, 
{17'b11111111110011001, 17'b00000000000001001, 17'b11111111111111111, 17'b00000000000101100, 17'b00000000000010001}, 
{17'b11111111111111111, 17'b00000000001001000, 17'b11111111110011011, 17'b00000000000101001, 17'b00000000000100010}, 
{17'b00000000000101001, 17'b11111111111010100, 17'b00000000000000000, 17'b11111111110001001, 17'b11111111111000000}, 
{17'b11111111111111111, 17'b11111111110111011, 17'b00000000000101101, 17'b00000000001101110, 17'b00000000000000000}, 
{17'b11111111111011110, 17'b11111111111011010, 17'b00000000000000000, 17'b00000000010010100, 17'b11111111110111011}, 
{17'b00000000000101011, 17'b00000000000111010, 17'b11111111110101000, 17'b11111111111111000, 17'b00000000000011111}, 
{17'b00000000000000000, 17'b00000000000101010, 17'b00000000000000010, 17'b11111111111001010, 17'b11111111101100000}, 
{17'b00000000000101101, 17'b00000000000010000, 17'b00000000001101011, 17'b11111111111101110, 17'b11111111110010010}, 
{17'b00000000000010111, 17'b11111111111110011, 17'b11111111110100011, 17'b11111111111110111, 17'b00000000010001001}, 
{17'b11111111110000110, 17'b11111111111000001, 17'b11111111111000111, 17'b00000000001100110, 17'b00000000000001000}, 
{17'b00000000001011000, 17'b11111111111010100, 17'b11111111111011101, 17'b11111111111000110, 17'b11111111111110000}, 
{17'b00000000000110001, 17'b11111111111110101, 17'b11111111110010110, 17'b11111111111111000, 17'b00000000000010010}, 
{17'b00000000001000010, 17'b00000000000001010, 17'b11111111111001000, 17'b00000000000000000, 17'b11111111110011111}, 
{17'b00000000000111011, 17'b11111111111101001, 17'b11111111111001001, 17'b00000000000110101, 17'b00000000000011000}, 
{17'b00000000000010001, 17'b11111111111111000, 17'b00000000001001100, 17'b11111111110010001, 17'b11111111111111010}, 
{17'b00000000000000000, 17'b00000000000011110, 17'b00000000001111100, 17'b11111111101111011, 17'b11111111101100001}, 
{17'b11111111111100110, 17'b00000000000011100, 17'b00000000000101101, 17'b11111111110100100, 17'b00000000010000101}, 
{17'b11111111111111111, 17'b00000000000101010, 17'b00000000001001000, 17'b00000000000001001, 17'b11111111101101101}, 
{17'b11111111111010100, 17'b00000000001011101, 17'b11111111111000110, 17'b00000000000000001, 17'b00000000001100011}, 
{17'b00000000000000110, 17'b00000000001000100, 17'b00000000000000111, 17'b11111111101000000, 17'b00000000010001100}, 
{17'b11111111110001010, 17'b11111111111000001, 17'b00000000000110110, 17'b00000000000111110, 17'b00000000000110011}, 
{17'b00000000000000001, 17'b00000000000111101, 17'b11111111111110110, 17'b11111111111011001, 17'b00000000000001000}, 
{17'b11111111111100101, 17'b00000000000111111, 17'b11111111101111111, 17'b00000000000100011, 17'b11111111111010111}, 
{17'b11111111111111011, 17'b00000000000100100, 17'b11111111111010100, 17'b11111111110011001, 17'b00000000010010111}, 
{17'b00000000001110010, 17'b00000000000010001, 17'b00000000001010011, 17'b11111111101101001, 17'b11111111110101111}, 
{17'b11111111111110000, 17'b11111111110011101, 17'b00000000001011101, 17'b00000000000010010, 17'b00000000000100000}
};

localparam logic signed [16:0] bias [5] = '{
17'b11111111111110000,  // -0.06223141402006149
17'b11111111111101111,  // -0.06270556896924973
17'b11111111111101110,  // -0.07014333456754684
17'b00000000000010101,  // 0.0820775106549263
17'b00000000000110111   // 0.2155742198228836
};
endpackage