// Width: 12
// NFRAC: 6
package dense_3_12_6;

localparam logic signed [11:0] weights [32][32] = '{ 
{12'b111111111100, 12'b111111100100, 12'b111111100110, 12'b111111110011, 12'b000000010101, 12'b000000000010, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b000000001000, 12'b111111011110, 12'b111111111100, 12'b000000110110, 12'b111111110000, 12'b111111000100, 12'b111111111101, 12'b000000000111, 12'b000000011011, 12'b111111101001, 12'b111110111011, 12'b111111111101, 12'b000000000011, 12'b111111100110, 12'b000000000000, 12'b000001000000, 12'b111110100010, 12'b111111110001, 12'b111111100111, 12'b111111110110, 12'b000000011011, 12'b111111110101}, 
{12'b000000101111, 12'b000001101110, 12'b000000011001, 12'b111111010101, 12'b000000001111, 12'b111111101110, 12'b111111111001, 12'b000001000101, 12'b000000000000, 12'b111111111111, 12'b111111111101, 12'b111111011010, 12'b111111110011, 12'b000000100010, 12'b111101111001, 12'b111111100001, 12'b111111111111, 12'b111111111111, 12'b111111111100, 12'b111111110101, 12'b111111101111, 12'b111111101110, 12'b000000000001, 12'b111111111111, 12'b111111111111, 12'b111110111011, 12'b000000000000, 12'b000000011110, 12'b111111111011, 12'b111111010011, 12'b000000000000, 12'b000000000010}, 
{12'b111111000000, 12'b000000001011, 12'b000000000000, 12'b000000010100, 12'b111111010111, 12'b000000000000, 12'b000000000000, 12'b111111001010, 12'b000000100010, 12'b111111101111, 12'b111111101111, 12'b111110100000, 12'b111111101100, 12'b000000100000, 12'b000000010000, 12'b111111111111, 12'b111111111000, 12'b111111111110, 12'b111111001011, 12'b000000000000, 12'b000000000111, 12'b000000000100, 12'b000000001101, 12'b000000111000, 12'b000000000010, 12'b111111001101, 12'b000000110001, 12'b000000000000, 12'b000000001010, 12'b111111111110, 12'b000000000000, 12'b000010010001}, 
{12'b000000110101, 12'b111111111111, 12'b111111110011, 12'b000001010011, 12'b000001001110, 12'b000000000000, 12'b000000000100, 12'b000000110100, 12'b111111100110, 12'b111111111111, 12'b111111001011, 12'b000000000111, 12'b000000010001, 12'b111111010000, 12'b000000000101, 12'b111111110101, 12'b111111111111, 12'b111111101000, 12'b000000000010, 12'b000000000011, 12'b000000000001, 12'b111111111011, 12'b000001001100, 12'b000000101011, 12'b000000101010, 12'b000000011111, 12'b000000101011, 12'b000000000000, 12'b111111111000, 12'b000000111001, 12'b000000011111, 12'b111111110100}, 
{12'b000001000000, 12'b111111111010, 12'b111111010011, 12'b111110011111, 12'b000000111101, 12'b000000000000, 12'b111111001011, 12'b111111011011, 12'b111111111010, 12'b111110011000, 12'b111101110010, 12'b000000111100, 12'b000001010101, 12'b000001000010, 12'b111110110110, 12'b111110011100, 12'b000000000000, 12'b111111101101, 12'b000000011001, 12'b000000010001, 12'b111111100111, 12'b111111111111, 12'b000001011100, 12'b111101010000, 12'b000000001011, 12'b111110101011, 12'b000000001000, 12'b111111100000, 12'b111111011001, 12'b111111111111, 12'b000000001000, 12'b000001001010}, 
{12'b000000000101, 12'b111111111010, 12'b111111011000, 12'b111111011110, 12'b000000101111, 12'b000000000000, 12'b111111011100, 12'b111111101110, 12'b111111001001, 12'b111111110111, 12'b111111111111, 12'b000000010100, 12'b000000000000, 12'b000000101101, 12'b111110111111, 12'b111111101111, 12'b000000001011, 12'b111111011010, 12'b111111100110, 12'b111111111111, 12'b000000000001, 12'b000000100110, 12'b000000111011, 12'b111111111110, 12'b111111111111, 12'b000000110011, 12'b111110111001, 12'b111111111111, 12'b111111100001, 12'b111111111011, 12'b111111111111, 12'b000000000000}, 
{12'b000000001000, 12'b111111010101, 12'b000000001101, 12'b111111111011, 12'b111111111111, 12'b000000010011, 12'b111111110010, 12'b111110101001, 12'b111111111111, 12'b111111100101, 12'b111111000101, 12'b000000111100, 12'b000000000000, 12'b000001010111, 12'b000001101010, 12'b000000000000, 12'b111111111111, 12'b111111010111, 12'b111111111000, 12'b000000100010, 12'b111110011111, 12'b000000010011, 12'b000000101001, 12'b000000000010, 12'b000000010011, 12'b000010011111, 12'b111111001101, 12'b111111110100, 12'b111111100111, 12'b000000111110, 12'b111111111001, 12'b111111101010}, 
{12'b111110110011, 12'b000000000011, 12'b111110101111, 12'b000000110111, 12'b000010000011, 12'b000000001110, 12'b000000000000, 12'b000000000110, 12'b111111111111, 12'b000000010000, 12'b000010100110, 12'b111111111111, 12'b000000110000, 12'b000001001111, 12'b000001100010, 12'b000010000110, 12'b000000000000, 12'b111111000010, 12'b000000101011, 12'b111111111111, 12'b111110101110, 12'b111111100010, 12'b000000000001, 12'b111111110101, 12'b111110111111, 12'b000011110000, 12'b111111100011, 12'b000000000000, 12'b000000000000, 12'b000001110001, 12'b000000001011, 12'b000000110010}, 
{12'b000000110110, 12'b111111111101, 12'b000000000000, 12'b111111111010, 12'b000000001010, 12'b111111111011, 12'b111111111111, 12'b000000010100, 12'b000000011011, 12'b111111011100, 12'b000000010001, 12'b000000010111, 12'b000000000001, 12'b000000101010, 12'b111111100011, 12'b111110011001, 12'b000000000000, 12'b111111111110, 12'b111111111100, 12'b111111000000, 12'b111111111111, 12'b000000000000, 12'b111111100110, 12'b111111111110, 12'b111111110011, 12'b000000010011, 12'b000000101111, 12'b111111110000, 12'b111111111001, 12'b111111111010, 12'b000000000011, 12'b111111001101}, 
{12'b111111101001, 12'b000000110001, 12'b000000000000, 12'b000000000000, 12'b000001100101, 12'b000000101001, 12'b111111111111, 12'b111110111000, 12'b000000001111, 12'b111110100110, 12'b111101001100, 12'b111111111111, 12'b000000000000, 12'b000000110110, 12'b000000001110, 12'b000000000000, 12'b111111010101, 12'b000000000000, 12'b000000000000, 12'b000000000111, 12'b000000011111, 12'b111111111100, 12'b111111010001, 12'b000000000001, 12'b111111111110, 12'b000010001010, 12'b000000101001, 12'b111111111111, 12'b111111110110, 12'b000001010101, 12'b111111111010, 12'b111111110100}, 
{12'b111110111101, 12'b000000010110, 12'b111111111011, 12'b111111111111, 12'b111111100000, 12'b111111001111, 12'b000000000110, 12'b000000010010, 12'b111111111111, 12'b111111101010, 12'b111110110110, 12'b000000011001, 12'b000000100110, 12'b000000000000, 12'b000001101011, 12'b111110111000, 12'b000000001101, 12'b111111001101, 12'b000000100100, 12'b111111111111, 12'b111111111011, 12'b000000001000, 12'b000000001111, 12'b000000000000, 12'b111111000000, 12'b000000000011, 12'b111110111000, 12'b111111111010, 12'b111111111111, 12'b000001010110, 12'b111111100111, 12'b000000000000}, 
{12'b111111111111, 12'b000000001110, 12'b000000000000, 12'b000000110010, 12'b111111110001, 12'b111111111010, 12'b000000000111, 12'b111111111111, 12'b111111111010, 12'b000001010010, 12'b000001011001, 12'b000000000000, 12'b111111010101, 12'b111110100110, 12'b111111111001, 12'b000000000000, 12'b000000000000, 12'b111111110111, 12'b111111000011, 12'b000000110000, 12'b000000000000, 12'b000000101111, 12'b111111111111, 12'b000001000111, 12'b000000001111, 12'b000000100111, 12'b000000111010, 12'b111111111001, 12'b111111001101, 12'b111111000111, 12'b111111111111, 12'b111110101010}, 
{12'b111111100011, 12'b111111111111, 12'b000000001111, 12'b111111001010, 12'b000000001011, 12'b111111111111, 12'b111111100100, 12'b111111111110, 12'b111111101111, 12'b000000000100, 12'b000000001001, 12'b111111110110, 12'b000000000010, 12'b000000011000, 12'b111110101111, 12'b111111100000, 12'b000000011101, 12'b111111101001, 12'b000000000000, 12'b111111111100, 12'b000000011000, 12'b000000000001, 12'b111111111100, 12'b000000000101, 12'b000000100010, 12'b111111110010, 12'b000000000000, 12'b111111000110, 12'b111111100110, 12'b111111111111, 12'b000000010110, 12'b000000000000}, 
{12'b111110111101, 12'b000000110101, 12'b111111111111, 12'b111111111111, 12'b111111111110, 12'b000000010110, 12'b111111111111, 12'b000001100010, 12'b111111111110, 12'b111111111111, 12'b000000011010, 12'b000000000101, 12'b000000000000, 12'b000000000000, 12'b000000001111, 12'b000000101010, 12'b000000010110, 12'b000000010101, 12'b111111111110, 12'b000000100111, 12'b000000001100, 12'b000000000101, 12'b111111111110, 12'b000000100000, 12'b111111110011, 12'b111111010100, 12'b111111110100, 12'b111111111111, 12'b000000001101, 12'b000000000011, 12'b000000011001, 12'b000000111101}, 
{12'b111111111101, 12'b111111001110, 12'b000000000110, 12'b111111111111, 12'b000001110101, 12'b111111100101, 12'b111110110110, 12'b000000000000, 12'b000000000000, 12'b111111111100, 12'b000000000110, 12'b000000110111, 12'b000000101001, 12'b000000000001, 12'b000000000100, 12'b111111101001, 12'b000000000100, 12'b111111111011, 12'b000000000000, 12'b000000001001, 12'b111111111011, 12'b000000000010, 12'b000000100010, 12'b000000000100, 12'b111111111110, 12'b111111001011, 12'b000000011010, 12'b111111111111, 12'b111111111111, 12'b111111110010, 12'b111111111101, 12'b111111110111}, 
{12'b000000000000, 12'b111111110111, 12'b111111101111, 12'b111111100100, 12'b111110111010, 12'b000001001110, 12'b000000000000, 12'b000000010101, 12'b000000100100, 12'b000000000001, 12'b111111111011, 12'b000000111100, 12'b000000011100, 12'b111111010001, 12'b111111101011, 12'b111111111010, 12'b111111001101, 12'b111111111101, 12'b000000000000, 12'b111111111111, 12'b000000010011, 12'b111111101110, 12'b000000000000, 12'b000000001001, 12'b111111111111, 12'b111111010100, 12'b000000010100, 12'b000000000000, 12'b000000000101, 12'b000000000001, 12'b111111010111, 12'b000000000010}, 
{12'b111111100110, 12'b111111101011, 12'b000000001001, 12'b111111110000, 12'b111111110100, 12'b000000001110, 12'b111111111111, 12'b000000000100, 12'b000000010000, 12'b111111111111, 12'b000000001111, 12'b111111101111, 12'b111111111110, 12'b111111111111, 12'b000000001101, 12'b111111111111, 12'b000000111110, 12'b111111111101, 12'b000000011111, 12'b111111101010, 12'b000000010100, 12'b000000001000, 12'b000000001010, 12'b000000000100, 12'b111111110101, 12'b111111011100, 12'b111111011110, 12'b000000001101, 12'b111111110101, 12'b000000000000, 12'b111111111100, 12'b000000011101}, 
{12'b111111111111, 12'b111111001100, 12'b111111001101, 12'b111111111111, 12'b000001010000, 12'b111111110100, 12'b000000000000, 12'b000000111101, 12'b111111101101, 12'b000000000000, 12'b111111001010, 12'b111111000001, 12'b000000111001, 12'b000000010011, 12'b111111110000, 12'b111111011100, 12'b000000010110, 12'b000000000000, 12'b111111100001, 12'b000000000011, 12'b000000001000, 12'b111111110100, 12'b000000100100, 12'b111110000010, 12'b000000000101, 12'b000000011110, 12'b111111111010, 12'b000000000001, 12'b111111100010, 12'b111111111111, 12'b111111100110, 12'b111111111100}, 
{12'b000000011011, 12'b000000101100, 12'b000001000110, 12'b111111100101, 12'b000000110101, 12'b000000100111, 12'b000000000000, 12'b000000111010, 12'b000000101101, 12'b111111110010, 12'b000001011001, 12'b111111010011, 12'b000001001111, 12'b000000111001, 12'b111101110110, 12'b111111111111, 12'b000000000000, 12'b000000000000, 12'b000000100001, 12'b111110111111, 12'b000000011100, 12'b111111100100, 12'b111111000001, 12'b111111101011, 12'b000000101010, 12'b111110101011, 12'b111111010101, 12'b111111111010, 12'b111111111111, 12'b111110110111, 12'b000000110010, 12'b000000000000}, 
{12'b111111111001, 12'b000000000000, 12'b111111111111, 12'b111111111111, 12'b111111010011, 12'b000000000001, 12'b000000000001, 12'b111111111110, 12'b111111111100, 12'b111111111010, 12'b000000010001, 12'b111111111111, 12'b000000001010, 12'b111111010100, 12'b000000001101, 12'b111111111111, 12'b000000010010, 12'b000000111001, 12'b111111010010, 12'b000000000110, 12'b111111110011, 12'b000000010000, 12'b000000011000, 12'b111111110101, 12'b111111011111, 12'b000000000010, 12'b000001101010, 12'b111111111100, 12'b111111111110, 12'b000000101001, 12'b000000000000, 12'b000001101110}, 
{12'b111110111101, 12'b000000000100, 12'b111111100100, 12'b000000110001, 12'b000000001110, 12'b111111111011, 12'b111111111111, 12'b111111111111, 12'b111111011001, 12'b111111111011, 12'b000000000000, 12'b111110111000, 12'b000000000001, 12'b111111111010, 12'b111111111111, 12'b111111111111, 12'b111111110001, 12'b000000000000, 12'b000000000000, 12'b000000010100, 12'b000000000010, 12'b000000000000, 12'b000000000000, 12'b111111111110, 12'b000000000000, 12'b000000000010, 12'b000001001010, 12'b111111111111, 12'b111111111111, 12'b111111111010, 12'b000000010110, 12'b111111111100}, 
{12'b111111111111, 12'b111111101100, 12'b000000011010, 12'b000000000101, 12'b111111010000, 12'b000000000000, 12'b000000100100, 12'b111111111111, 12'b000000000000, 12'b111111110011, 12'b000000001110, 12'b000000000010, 12'b000000101001, 12'b111110111001, 12'b111111110011, 12'b111111111101, 12'b000000011011, 12'b111111001110, 12'b000000000010, 12'b111110011111, 12'b111111111101, 12'b111111110000, 12'b111111111010, 12'b000000100101, 12'b111111110110, 12'b111111011100, 12'b000000001011, 12'b000000000000, 12'b000000110010, 12'b000001000010, 12'b111111010110, 12'b111111000110}, 
{12'b000000001000, 12'b000000000011, 12'b111111001010, 12'b111111111000, 12'b111111111111, 12'b000000000000, 12'b000000001101, 12'b000000110100, 12'b000000000000, 12'b000000000010, 12'b000000001000, 12'b111110111010, 12'b111111110111, 12'b111110110010, 12'b000000111101, 12'b000000000000, 12'b111111111111, 12'b111110101101, 12'b111111111111, 12'b111111110110, 12'b111111111101, 12'b000000000000, 12'b000000000111, 12'b111111101100, 12'b000000000110, 12'b000000110100, 12'b000000110110, 12'b000000110001, 12'b000000100111, 12'b000000000000, 12'b000000001110, 12'b000001100100}, 
{12'b111111111100, 12'b111111100001, 12'b000000110001, 12'b111111110010, 12'b000000001000, 12'b000000010101, 12'b111111111111, 12'b111111011011, 12'b111111110101, 12'b111110110011, 12'b000000111001, 12'b000000000000, 12'b000000110101, 12'b000001010101, 12'b111111110001, 12'b111110010000, 12'b111111110010, 12'b000000111100, 12'b111111011011, 12'b111111100101, 12'b000000000111, 12'b000000000000, 12'b111110111010, 12'b111111100111, 12'b111111111010, 12'b111111110000, 12'b000000001110, 12'b000001011010, 12'b000000011111, 12'b111111111111, 12'b000000001010, 12'b000000000011}, 
{12'b000000000101, 12'b000000111010, 12'b000000000000, 12'b000000100101, 12'b000001101010, 12'b111111101010, 12'b111111111111, 12'b111111111010, 12'b000000100101, 12'b111111100111, 12'b111111111111, 12'b000000101010, 12'b000000000001, 12'b000000000011, 12'b111100111100, 12'b111111110101, 12'b000000000000, 12'b000000011001, 12'b111111111111, 12'b000000100110, 12'b111111111111, 12'b111111101001, 12'b111110111000, 12'b000000010000, 12'b000000100100, 12'b111101110010, 12'b111111111111, 12'b000000000000, 12'b000001000101, 12'b111110011001, 12'b000000000000, 12'b111111111111}, 
{12'b000000000001, 12'b111111010100, 12'b000000000110, 12'b111111111110, 12'b000000000110, 12'b000001000011, 12'b111110100011, 12'b000000000100, 12'b000000110110, 12'b111111010100, 12'b111111111101, 12'b000000000110, 12'b111111111110, 12'b000000010110, 12'b000000001101, 12'b111111111101, 12'b000000001000, 12'b000000000000, 12'b000000000010, 12'b000000110000, 12'b111111111100, 12'b111111000010, 12'b111110110010, 12'b111111100111, 12'b111110110100, 12'b000000011010, 12'b000001001111, 12'b000000101111, 12'b111111111110, 12'b111111010000, 12'b111111011000, 12'b000000000111}, 
{12'b000000000110, 12'b111111000010, 12'b111111111101, 12'b000000010011, 12'b111111000010, 12'b000000010101, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b000000000000, 12'b000000100001, 12'b111111111101, 12'b000000000001, 12'b000000000000, 12'b000000010000, 12'b111111111101, 12'b000000000000, 12'b111111111111, 12'b111111010110, 12'b111110111111, 12'b111111111111, 12'b111110111011, 12'b111111011001, 12'b111111010000, 12'b000001110001, 12'b000000000010, 12'b111111111010, 12'b000000101000, 12'b000001110010, 12'b000000110010, 12'b111101111000, 12'b111111101000}, 
{12'b000000110000, 12'b111111111111, 12'b000000100000, 12'b111111111101, 12'b000000111101, 12'b111111101101, 12'b000000001001, 12'b000000110101, 12'b000000100010, 12'b111110111101, 12'b111111111000, 12'b000000001111, 12'b000000001000, 12'b111111111110, 12'b000000001010, 12'b000000000000, 12'b000000101110, 12'b000000000100, 12'b000000101111, 12'b111111110111, 12'b111111101111, 12'b111111110110, 12'b111111111111, 12'b000000100110, 12'b111111100110, 12'b111111111111, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000100101, 12'b111111010110, 12'b111111111101}, 
{12'b111111111111, 12'b111111111100, 12'b111111000100, 12'b000000100100, 12'b000000011100, 12'b111111110001, 12'b111111111111, 12'b111111100010, 12'b000000000000, 12'b111111111111, 12'b111111011001, 12'b111111100000, 12'b000000111101, 12'b000000000000, 12'b111111101111, 12'b111111111111, 12'b000000011011, 12'b111111111111, 12'b111111111111, 12'b111111100100, 12'b000000101000, 12'b000000000000, 12'b000000010011, 12'b111111111100, 12'b000000010100, 12'b000000000000, 12'b000000000000, 12'b000000011110, 12'b111111100111, 12'b111111111010, 12'b000000010100, 12'b111111110010}, 
{12'b111111111101, 12'b111111011000, 12'b000001001100, 12'b111111110111, 12'b000000011001, 12'b111111011011, 12'b000000000000, 12'b000000000100, 12'b111111000010, 12'b111111111110, 12'b111111110000, 12'b000000000111, 12'b111111010110, 12'b000000010001, 12'b000000011001, 12'b000000001110, 12'b000000001010, 12'b111111111011, 12'b111110100101, 12'b111111111110, 12'b111111111000, 12'b000000010001, 12'b111111110001, 12'b111111111111, 12'b000000011001, 12'b111111111010, 12'b111111111110, 12'b000000110001, 12'b111111001101, 12'b111111011010, 12'b000000101100, 12'b000000000100}, 
{12'b000000110111, 12'b000000011001, 12'b000000000000, 12'b111111101011, 12'b111111110101, 12'b111111111111, 12'b000000000000, 12'b111111110111, 12'b111111110000, 12'b111111110000, 12'b000000000000, 12'b000000010100, 12'b000000000000, 12'b000000000110, 12'b111111111010, 12'b000000000000, 12'b111111101100, 12'b000000000000, 12'b111111111101, 12'b111111111111, 12'b000000000000, 12'b000000000111, 12'b000000001100, 12'b000000000000, 12'b000000000000, 12'b111110110001, 12'b111111100110, 12'b000000000000, 12'b000000000010, 12'b000000000000, 12'b111111101001, 12'b000000000010}, 
{12'b000000011000, 12'b111101111010, 12'b111111111111, 12'b111111110110, 12'b111111100010, 12'b111111111110, 12'b000000000000, 12'b000001000110, 12'b111111111010, 12'b111111111101, 12'b000000001010, 12'b111110101011, 12'b000000000011, 12'b111111000111, 12'b000001011100, 12'b111111111001, 12'b111111100011, 12'b111110111001, 12'b111111111110, 12'b111110100101, 12'b111110011000, 12'b111111111111, 12'b000000000000, 12'b000000000000, 12'b000000011111, 12'b111111111110, 12'b111111011001, 12'b111111110110, 12'b111111111101, 12'b000000000000, 12'b111111111011, 12'b111110100110}
};

localparam logic signed [11:0] bias [32] = '{
12'b000000100001,  // 0.5280959606170654
12'b000000110101,  // 0.8414360880851746
12'b000000011001,  // 0.397830605506897
12'b000000011010,  // 0.4105983078479767
12'b111100010101,  // -3.657735586166382
12'b111111000110,  // -0.8977976441383362
12'b000001101101,  // 1.7051936388015747
12'b111110101110,  // -1.2765135765075684
12'b111111011010,  // -0.5837795734405518
12'b000010101100,  // 2.699671983718872
12'b000000001101,  // 0.2170683741569519
12'b000000111000,  // 0.8814588785171509
12'b111101010111,  // -2.634300947189331
12'b111110000111,  // -1.877297282218933
12'b000001101010,  // 1.6625694036483765
12'b000010101111,  // 2.7459704875946045
12'b111111100001,  // -0.47838035225868225
12'b000001101100,  // 1.6984987258911133
12'b000000110110,  // 0.8548859357833862
12'b000001000000,  // 1.0045719146728516
12'b000001011010,  // 1.4197649955749512
12'b000000110101,  // 0.832463800907135
12'b000000100010,  // 0.5434179306030273
12'b000000111011,  // 0.9277304410934448
12'b111111101010,  // -0.3426123857498169
12'b111111011100,  // -0.5587119460105896
12'b111111011000,  // -0.6208624839782715
12'b111110101110,  // -1.2802538871765137
12'b000000000011,  // 0.05940237268805504
12'b111111001011,  // -0.8213341236114502
12'b000000111000,  // 0.8783953189849854
12'b111111000011   // -0.949700653553009
};
endpackage