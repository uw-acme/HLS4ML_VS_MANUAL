// Width: 16
// NFRAC: 10
package dense_3_16_10;

localparam logic signed [15:0] weights [32][32] = '{ 
{16'b1111111111001101, 16'b1111111001000000, 16'b1111111001100000, 16'b1111111100111100, 16'b0000000101011111, 16'b0000000000101100, 16'b1111111111110010, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000010000001, 16'b1111110111100100, 16'b1111111111000010, 16'b0000001101100011, 16'b1111111100001000, 16'b1111110001000100, 16'b1111111111011010, 16'b0000000001110010, 16'b0000000110111101, 16'b1111111010011011, 16'b1111101110111100, 16'b1111111111010000, 16'b0000000000110010, 16'b1111111001100011, 16'b0000000000000000, 16'b0000010000001100, 16'b1111101000101100, 16'b1111111100011101, 16'b1111111001110010, 16'b1111111101100110, 16'b0000000110110001, 16'b1111111101011100}, 
{16'b0000001011111101, 16'b0000011011101011, 16'b0000000110011011, 16'b1111110101011110, 16'b0000000011111010, 16'b1111111011101000, 16'b1111111110010000, 16'b0000010001011100, 16'b0000000000000110, 16'b1111111111111111, 16'b1111111111011111, 16'b1111110110100101, 16'b1111111100110001, 16'b0000001000101001, 16'b1111011110010011, 16'b1111111000011101, 16'b1111111111111111, 16'b1111111111110111, 16'b1111111111001010, 16'b1111111101010111, 16'b1111111011110111, 16'b1111111011100110, 16'b0000000000010001, 16'b1111111111111110, 16'b1111111111111001, 16'b1111101110110110, 16'b0000000000001100, 16'b0000000111100010, 16'b1111111110111111, 16'b1111110100111101, 16'b0000000000000010, 16'b0000000000100110}, 
{16'b1111110000001111, 16'b0000000010111100, 16'b0000000000001010, 16'b0000000101001010, 16'b1111110101111010, 16'b0000000000000000, 16'b0000000000000001, 16'b1111110010100100, 16'b0000001000100100, 16'b1111111011110011, 16'b1111111011110110, 16'b1111101000001101, 16'b1111111011000001, 16'b0000001000001011, 16'b0000000100001110, 16'b1111111111111110, 16'b1111111110001010, 16'b1111111111100111, 16'b1111110010111101, 16'b0000000000000011, 16'b0000000001111111, 16'b0000000001000110, 16'b0000000011010110, 16'b0000001110000101, 16'b0000000000100110, 16'b1111110011011000, 16'b0000001100010001, 16'b0000000000000000, 16'b0000000010101001, 16'b1111111111101001, 16'b0000000000000000, 16'b0000100100010011}, 
{16'b0000001101011001, 16'b1111111111111111, 16'b1111111100111000, 16'b0000010100111100, 16'b0000010011101001, 16'b0000000000000000, 16'b0000000001001011, 16'b0000001101000001, 16'b1111111001101010, 16'b1111111111111111, 16'b1111110010110100, 16'b0000000001111010, 16'b0000000100010000, 16'b1111110100000010, 16'b0000000001011111, 16'b1111111101011100, 16'b1111111111111111, 16'b1111111010001011, 16'b0000000000100111, 16'b0000000000111000, 16'b0000000000010000, 16'b1111111110110101, 16'b0000010011000110, 16'b0000001010111110, 16'b0000001010100010, 16'b0000000111111100, 16'b0000001010111011, 16'b0000000000000000, 16'b1111111110000111, 16'b0000001110011111, 16'b0000000111111111, 16'b1111111101001100}, 
{16'b0000010000000000, 16'b1111111110100000, 16'b1111110100111010, 16'b1111100111111100, 16'b0000001111010001, 16'b0000000000000000, 16'b1111110010110111, 16'b1111110110111101, 16'b1111111110100000, 16'b1111100110000110, 16'b1111011100101001, 16'b0000001111001000, 16'b0000010101011001, 16'b0000010000101111, 16'b1111101101100110, 16'b1111100111001100, 16'b0000000000000000, 16'b1111111011011110, 16'b0000000110011011, 16'b0000000100011100, 16'b1111111001111110, 16'b1111111111110010, 16'b0000010111000101, 16'b1111010100000000, 16'b0000000010110100, 16'b1111101010111011, 16'b0000000010000110, 16'b1111111000000011, 16'b1111110110011100, 16'b1111111111111111, 16'b0000000010001111, 16'b0000010010100100}, 
{16'b0000000001011000, 16'b1111111110101011, 16'b1111110110001011, 16'b1111110111101010, 16'b0000001011111001, 16'b0000000000000000, 16'b1111110111000011, 16'b1111111011101001, 16'b1111110010010011, 16'b1111111101111100, 16'b1111111111111111, 16'b0000000101001000, 16'b0000000000000000, 16'b0000001011011100, 16'b1111101111110100, 16'b1111111011111010, 16'b0000000010110110, 16'b1111110110100111, 16'b1111111001101011, 16'b1111111111111111, 16'b0000000000011000, 16'b0000001001100101, 16'b0000001110111100, 16'b1111111111101010, 16'b1111111111111111, 16'b0000001100110100, 16'b1111101110011010, 16'b1111111111111111, 16'b1111111000011011, 16'b1111111110110100, 16'b1111111111111001, 16'b0000000000001101}, 
{16'b0000000010000101, 16'b1111110101010111, 16'b0000000011011101, 16'b1111111110110001, 16'b1111111111110000, 16'b0000000100110110, 16'b1111111100100110, 16'b1111101010010101, 16'b1111111111111111, 16'b1111111001010101, 16'b1111110001011000, 16'b0000001111000111, 16'b0000000000001110, 16'b0000010101111001, 16'b0000011010100001, 16'b0000000000000101, 16'b1111111111111111, 16'b1111110101111010, 16'b1111111110000001, 16'b0000001000101111, 16'b1111100111111111, 16'b0000000100111111, 16'b0000001010011100, 16'b0000000000100110, 16'b0000000100110011, 16'b0000100111110010, 16'b1111110011011000, 16'b1111111101000110, 16'b1111111001111011, 16'b0000001111100101, 16'b1111111110011011, 16'b1111111010100101}, 
{16'b1111101100111010, 16'b0000000000110000, 16'b1111101011110111, 16'b0000001101111011, 16'b0000100000111001, 16'b0000000011101101, 16'b0000000000000111, 16'b0000000001100000, 16'b1111111111111111, 16'b0000000100000110, 16'b0000101001101000, 16'b1111111111111111, 16'b0000001100001100, 16'b0000010011111011, 16'b0000011000100110, 16'b0000100001100110, 16'b0000000000000000, 16'b1111110000101100, 16'b0000001010110000, 16'b1111111111110100, 16'b1111101011100101, 16'b1111111000101111, 16'b0000000000011011, 16'b1111111101010110, 16'b1111101111111101, 16'b0000111100000001, 16'b1111111000111110, 16'b0000000000000000, 16'b0000000000000000, 16'b0000011100010000, 16'b0000000010110101, 16'b0000001100100010}, 
{16'b0000001101100000, 16'b1111111111011000, 16'b0000000000000000, 16'b1111111110100111, 16'b0000000010100111, 16'b1111111110110010, 16'b1111111111111111, 16'b0000000101000001, 16'b0000000110110000, 16'b1111110111001110, 16'b0000000100011110, 16'b0000000101111111, 16'b0000000000011000, 16'b0000001010101001, 16'b1111111000110011, 16'b1111100110011111, 16'b0000000000000000, 16'b1111111111100011, 16'b1111111111001001, 16'b1111110000000010, 16'b1111111111111101, 16'b0000000000000000, 16'b1111111001100000, 16'b1111111111100011, 16'b1111111100111101, 16'b0000000100111111, 16'b0000001011111101, 16'b1111111100001011, 16'b1111111110011011, 16'b1111111110101101, 16'b0000000000110111, 16'b1111110011011100}, 
{16'b1111111010010100, 16'b0000001100010011, 16'b0000000000000000, 16'b0000000000000000, 16'b0000011001010110, 16'b0000001010010011, 16'b1111111111111111, 16'b1111101110001111, 16'b0000000011110001, 16'b1111101001101011, 16'b1111010011000110, 16'b1111111111111111, 16'b0000000000000000, 16'b0000001101101110, 16'b0000000011100011, 16'b0000000000000000, 16'b1111110101011111, 16'b0000000000000000, 16'b0000000000001101, 16'b0000000001111100, 16'b0000000111110011, 16'b1111111111001011, 16'b1111110100011110, 16'b0000000000010000, 16'b1111111111101000, 16'b0000100010100110, 16'b0000001010011100, 16'b1111111111111111, 16'b1111111101101110, 16'b0000010101011000, 16'b1111111110101110, 16'b1111111101001100}, 
{16'b1111101111010000, 16'b0000000101100110, 16'b1111111110111000, 16'b1111111111111111, 16'b1111111000000111, 16'b1111110011111010, 16'b0000000001100010, 16'b0000000100100111, 16'b1111111111111111, 16'b1111111010100001, 16'b1111101101101011, 16'b0000000110011011, 16'b0000001001101110, 16'b0000000000000000, 16'b0000011010110110, 16'b1111101110000001, 16'b0000000011010100, 16'b1111110011011111, 16'b0000001001000001, 16'b1111111111111111, 16'b1111111110110001, 16'b0000000010001111, 16'b0000000011111011, 16'b0000000000000000, 16'b1111110000001100, 16'b0000000000111111, 16'b1111101110000111, 16'b1111111110101110, 16'b1111111111111111, 16'b0000010101100111, 16'b1111111001111010, 16'b0000000000000000}, 
{16'b1111111111111111, 16'b0000000011101011, 16'b0000000000000000, 16'b0000001100100001, 16'b1111111100010000, 16'b1111111110100111, 16'b0000000001110111, 16'b1111111111110100, 16'b1111111110100001, 16'b0000010100100000, 16'b0000010110010111, 16'b0000000000000001, 16'b1111110101010110, 16'b1111101001100001, 16'b1111111110011000, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111101111101, 16'b1111110000110000, 16'b0000001100001111, 16'b0000000000000100, 16'b0000001011110111, 16'b1111111111111111, 16'b0000010001111111, 16'b0000000011111101, 16'b0000001001110011, 16'b0000001110100100, 16'b1111111110010110, 16'b1111110011011110, 16'b1111110001111001, 16'b1111111111110101, 16'b1111101010100110}, 
{16'b1111111000110000, 16'b1111111111111111, 16'b0000000011110100, 16'b1111110010100110, 16'b0000000010110000, 16'b1111111111111111, 16'b1111111001000011, 16'b1111111111101100, 16'b1111111011111111, 16'b0000000001001100, 16'b0000000010011111, 16'b1111111101101101, 16'b0000000000100001, 16'b0000000110000000, 16'b1111101011111111, 16'b1111111000001010, 16'b0000000111010011, 16'b1111111010010101, 16'b0000000000000000, 16'b1111111111001100, 16'b0000000110001011, 16'b0000000000010000, 16'b1111111111000000, 16'b0000000001010111, 16'b0000001000100111, 16'b1111111100101011, 16'b0000000000000000, 16'b1111110001100010, 16'b1111111001101111, 16'b1111111111110001, 16'b0000000101100011, 16'b0000000000000000}, 
{16'b1111101111010111, 16'b0000001101011100, 16'b1111111111111111, 16'b1111111111110010, 16'b1111111111101100, 16'b0000000101100111, 16'b1111111111111111, 16'b0000011000101101, 16'b1111111111100001, 16'b1111111111111111, 16'b0000000110100101, 16'b0000000001010011, 16'b0000000000001101, 16'b0000000000000000, 16'b0000000011111001, 16'b0000001010100100, 16'b0000000101101100, 16'b0000000101010101, 16'b1111111111101110, 16'b0000001001110101, 16'b0000000011001110, 16'b0000000001010010, 16'b1111111111101110, 16'b0000001000001000, 16'b1111111100110100, 16'b1111110101001001, 16'b1111111101000010, 16'b1111111111111111, 16'b0000000011010000, 16'b0000000000111100, 16'b0000000110010000, 16'b0000001111010101}, 
{16'b1111111111011001, 16'b1111110011100010, 16'b0000000001101001, 16'b1111111111111110, 16'b0000011101010100, 16'b1111111001010111, 16'b1111101101101101, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111001011, 16'b0000000001100011, 16'b0000001101111110, 16'b0000001010010011, 16'b0000000000010101, 16'b0000000001000100, 16'b1111111010011010, 16'b0000000001000100, 16'b1111111110110010, 16'b0000000000000000, 16'b0000000010011010, 16'b1111111110110011, 16'b0000000000100111, 16'b0000001000100001, 16'b0000000001001011, 16'b1111111111100111, 16'b1111110010110010, 16'b0000000110100000, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111100100110, 16'b1111111111010100, 16'b1111111101111111}, 
{16'b0000000000001110, 16'b1111111101111110, 16'b1111111011111101, 16'b1111111001000000, 16'b1111101110100000, 16'b0000010011100000, 16'b0000000000000000, 16'b0000000101011001, 16'b0000001001001011, 16'b0000000000011010, 16'b1111111110111010, 16'b0000001111001110, 16'b0000000111001010, 16'b1111110100010011, 16'b1111111010110011, 16'b1111111110101011, 16'b1111110011010000, 16'b1111111111011100, 16'b0000000000000000, 16'b1111111111110110, 16'b0000000100111111, 16'b1111111011100111, 16'b0000000000000000, 16'b0000000010011101, 16'b1111111111111111, 16'b1111110101000100, 16'b0000000101000000, 16'b0000000000000000, 16'b0000000001011011, 16'b0000000000010110, 16'b1111110101111000, 16'b0000000000101010}, 
{16'b1111111001101110, 16'b1111111010111101, 16'b0000000010011100, 16'b1111111100000001, 16'b1111111101001000, 16'b0000000011101101, 16'b1111111111110101, 16'b0000000001000111, 16'b0000000100001100, 16'b1111111111111111, 16'b0000000011111101, 16'b1111111011111011, 16'b1111111111101100, 16'b1111111111111111, 16'b0000000011010011, 16'b1111111111111111, 16'b0000001111101000, 16'b1111111111011100, 16'b0000000111111100, 16'b1111111010100100, 16'b0000000101000100, 16'b0000000010000000, 16'b0000000010101100, 16'b0000000001001010, 16'b1111111101011001, 16'b1111110111000101, 16'b1111110111101101, 16'b0000000011011101, 16'b1111111101010100, 16'b0000000000000001, 16'b1111111111000111, 16'b0000000111011011}, 
{16'b1111111111111111, 16'b1111110011000010, 16'b1111110011010011, 16'b1111111111111111, 16'b0000010100001100, 16'b1111111101000110, 16'b0000000000000000, 16'b0000001111011101, 16'b1111111011010001, 16'b0000000000000000, 16'b1111110010101000, 16'b1111110000010100, 16'b0000001110010110, 16'b0000000100110101, 16'b1111111100000111, 16'b1111110111001111, 16'b0000000101100001, 16'b0000000000000000, 16'b1111111000011001, 16'b0000000000110110, 16'b0000000010001110, 16'b1111111101001010, 16'b0000001001000101, 16'b1111100000101001, 16'b0000000001010011, 16'b0000000111101001, 16'b1111111110101011, 16'b0000000000011110, 16'b1111111000100010, 16'b1111111111111111, 16'b1111111001100100, 16'b1111111111001110}, 
{16'b0000000110110011, 16'b0000001011000010, 16'b0000010001100111, 16'b1111111001011101, 16'b0000001101010100, 16'b0000001001110011, 16'b0000000000000001, 16'b0000001110100100, 16'b0000001011011011, 16'b1111111100100101, 16'b0000010110011100, 16'b1111110100110100, 16'b0000010011111000, 16'b0000001110010010, 16'b1111011101101010, 16'b1111111111111110, 16'b0000000000000000, 16'b0000000000001011, 16'b0000001000010100, 16'b1111101111111001, 16'b0000000111000101, 16'b1111111001001101, 16'b1111110000010011, 16'b1111111010111110, 16'b0000001010100010, 16'b1111101010111000, 16'b1111110101011100, 16'b1111111110101011, 16'b1111111111111111, 16'b1111101101111100, 16'b0000001100101001, 16'b0000000000000000}, 
{16'b1111111110011011, 16'b0000000000000001, 16'b1111111111111111, 16'b1111111111111111, 16'b1111110100110000, 16'b0000000000010010, 16'b0000000000010000, 16'b1111111111100001, 16'b1111111111001110, 16'b1111111110100001, 16'b0000000100011100, 16'b1111111111111110, 16'b0000000010101001, 16'b1111110101000011, 16'b0000000011011010, 16'b1111111111111110, 16'b0000000100100000, 16'b0000001110010100, 16'b1111110100101101, 16'b0000000001101010, 16'b1111111100110101, 16'b0000000100000111, 16'b0000000110000101, 16'b1111111101010001, 16'b1111110111111101, 16'b0000000000101010, 16'b0000011010100010, 16'b1111111111001110, 16'b1111111111100000, 16'b0000001010011000, 16'b0000000000000000, 16'b0000011011100101}, 
{16'b1111101111010011, 16'b0000000001001010, 16'b1111111001000100, 16'b0000001100010000, 16'b0000000011100000, 16'b1111111110111111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111110110010011, 16'b1111111110111100, 16'b0000000000000000, 16'b1111101110001110, 16'b0000000000011001, 16'b1111111110101110, 16'b1111111111111010, 16'b1111111111111111, 16'b1111111100010001, 16'b0000000000001011, 16'b0000000000000110, 16'b0000000101000100, 16'b0000000000100011, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111101111, 16'b0000000000000000, 16'b0000000000100101, 16'b0000010010100110, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111110101100, 16'b0000000101100110, 16'b1111111111001011}, 
{16'b1111111111111100, 16'b1111111011001010, 16'b0000000110100010, 16'b0000000001010001, 16'b1111110100000110, 16'b0000000000000001, 16'b0000001001001001, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111100110110, 16'b0000000011101011, 16'b0000000000100110, 16'b0000001010010110, 16'b1111101110011101, 16'b1111111100111110, 16'b1111111111011100, 16'b0000000110111010, 16'b1111110011101101, 16'b0000000000101011, 16'b1111100111110110, 16'b1111111111011001, 16'b1111111100001100, 16'b1111111110101101, 16'b0000001001011101, 16'b1111111101100111, 16'b1111110111000000, 16'b0000000010111001, 16'b0000000000000000, 16'b0000001100101010, 16'b0000010000101111, 16'b1111110101100000, 16'b1111110001101000}, 
{16'b0000000010001010, 16'b0000000000110100, 16'b1111110010101111, 16'b1111111110001011, 16'b1111111111111111, 16'b0000000000000100, 16'b0000000011011001, 16'b0000001101001010, 16'b0000000000000000, 16'b0000000000101001, 16'b0000000010001111, 16'b1111101110101111, 16'b1111111101110111, 16'b1111101100101011, 16'b0000001111011000, 16'b0000000000000000, 16'b1111111111111110, 16'b1111101011011111, 16'b1111111111111111, 16'b1111111101100111, 16'b1111111111010101, 16'b0000000000000000, 16'b0000000001111111, 16'b1111111011001100, 16'b0000000001101100, 16'b0000001101001001, 16'b0000001101101001, 16'b0000001100011111, 16'b0000001001110110, 16'b0000000000000000, 16'b0000000011101001, 16'b0000011001000100}, 
{16'b1111111111001100, 16'b1111111000011000, 16'b0000001100011101, 16'b1111111100101101, 16'b0000000010001110, 16'b0000000101010111, 16'b1111111111111111, 16'b1111110110110100, 16'b1111111101010001, 16'b1111101100110001, 16'b0000001110010100, 16'b0000000000000111, 16'b0000001101011010, 16'b0000010101011100, 16'b1111111100010001, 16'b1111100100001000, 16'b1111111100101011, 16'b0000001111000010, 16'b1111110110111100, 16'b1111111001010100, 16'b0000000001111001, 16'b0000000000000010, 16'b1111101110100011, 16'b1111111001111000, 16'b1111111110101111, 16'b1111111100000110, 16'b0000000011100101, 16'b0000010110100000, 16'b0000000111110110, 16'b1111111111111111, 16'b0000000010100101, 16'b0000000000111000}, 
{16'b0000000001010110, 16'b0000001110100001, 16'b0000000000000000, 16'b0000001001011101, 16'b0000011010100110, 16'b1111111010100010, 16'b1111111111111111, 16'b1111111110100101, 16'b0000001001011000, 16'b1111111001110111, 16'b1111111111111101, 16'b0000001010101010, 16'b0000000000010001, 16'b0000000000111000, 16'b1111001111001000, 16'b1111111101011101, 16'b0000000000000000, 16'b0000000110011011, 16'b1111111111111001, 16'b0000001001100011, 16'b1111111111111111, 16'b1111111010011110, 16'b1111101110000001, 16'b0000000100001011, 16'b0000001001001001, 16'b1111011100100000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000010001011010, 16'b1111100110010110, 16'b0000000000000011, 16'b1111111111110011}, 
{16'b0000000000010011, 16'b1111110101001000, 16'b0000000001101110, 16'b1111111111100001, 16'b0000000001101010, 16'b0000010000111011, 16'b1111101000110011, 16'b0000000001000110, 16'b0000001101100011, 16'b1111110101001101, 16'b1111111111010000, 16'b0000000001100100, 16'b1111111111101101, 16'b0000000101101110, 16'b0000000011011011, 16'b1111111111011101, 16'b0000000010001001, 16'b0000000000000000, 16'b0000000000101100, 16'b0000001100001001, 16'b1111111111000110, 16'b1111110000100000, 16'b1111101100101001, 16'b1111111001110011, 16'b1111101101000110, 16'b0000000110101010, 16'b0000010011111100, 16'b0000001011110011, 16'b1111111111101010, 16'b1111110100000100, 16'b1111110110000011, 16'b0000000001111010}, 
{16'b0000000001101010, 16'b1111110000101101, 16'b1111111111011101, 16'b0000000100110100, 16'b1111110000101100, 16'b0000000101011011, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b0000001000011101, 16'b1111111111011100, 16'b0000000000010011, 16'b0000000000000000, 16'b0000000100000100, 16'b1111111111011101, 16'b0000000000000101, 16'b1111111111111110, 16'b1111110101101100, 16'b1111101111110100, 16'b1111111111111110, 16'b1111101110111010, 16'b1111110110010111, 16'b1111110100000110, 16'b0000011100011111, 16'b0000000000100100, 16'b1111111110100001, 16'b0000001010001001, 16'b0000011100101110, 16'b0000001100101000, 16'b1111011110000100, 16'b1111111010000100}, 
{16'b0000001100000001, 16'b1111111111111111, 16'b0000001000000010, 16'b1111111111010111, 16'b0000001111011110, 16'b1111111011011011, 16'b0000000010010001, 16'b0000001101011000, 16'b0000001000100100, 16'b1111101111010010, 16'b1111111110000001, 16'b0000000011111011, 16'b0000000010001101, 16'b1111111111100010, 16'b0000000010101101, 16'b0000000000000000, 16'b0000001011100110, 16'b0000000001000111, 16'b0000001011111110, 16'b1111111101111001, 16'b1111111011111011, 16'b1111111101100110, 16'b1111111111111111, 16'b0000001001101010, 16'b1111111001100001, 16'b1111111111110011, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000001001010110, 16'b1111110101101111, 16'b1111111111010000}, 
{16'b1111111111111110, 16'b1111111111000000, 16'b1111110001000111, 16'b0000001001000110, 16'b0000000111001001, 16'b1111111100011111, 16'b1111111111111111, 16'b1111111000101111, 16'b0000000000001101, 16'b1111111111111111, 16'b1111110110010110, 16'b1111111000000111, 16'b0000001111010101, 16'b0000000000000000, 16'b1111111011111010, 16'b1111111111111111, 16'b0000000110110110, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111001000101, 16'b0000001010000111, 16'b0000000000000000, 16'b0000000100111111, 16'b1111111111000101, 16'b0000000101000001, 16'b0000000000000100, 16'b0000000000000000, 16'b0000000111101101, 16'b1111111001110110, 16'b1111111110100001, 16'b0000000101001000, 16'b1111111100100111}, 
{16'b1111111111011101, 16'b1111110110001000, 16'b0000010011000001, 16'b1111111101111010, 16'b0000000110010010, 16'b1111110110110110, 16'b0000000000000000, 16'b0000000001000110, 16'b1111110000101010, 16'b1111111111100101, 16'b1111111100000010, 16'b0000000001110111, 16'b1111110101100000, 16'b0000000100011010, 16'b0000000110011110, 16'b0000000011100000, 16'b0000000010101111, 16'b1111111110110010, 16'b1111101001010101, 16'b1111111111100100, 16'b1111111110001011, 16'b0000000100011110, 16'b1111111100011100, 16'b1111111111111111, 16'b0000000110010100, 16'b1111111110100010, 16'b1111111111100010, 16'b0000001100011100, 16'b1111110011010000, 16'b1111110110100011, 16'b0000001011001110, 16'b0000000001001001}, 
{16'b0000001101110010, 16'b0000000110011100, 16'b0000000000000001, 16'b1111111010111010, 16'b1111111101011111, 16'b1111111111111110, 16'b0000000000000000, 16'b1111111101110010, 16'b1111111100000001, 16'b1111111100001101, 16'b0000000000000000, 16'b0000000101000100, 16'b0000000000001101, 16'b0000000001101100, 16'b1111111110100100, 16'b0000000000001011, 16'b1111111011000101, 16'b0000000000000001, 16'b1111111111011011, 16'b1111111111111110, 16'b0000000000000100, 16'b0000000001111001, 16'b0000000011000111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111101100011101, 16'b1111111001100111, 16'b0000000000001101, 16'b0000000000101001, 16'b0000000000000010, 16'b1111111010010101, 16'b0000000000101011}, 
{16'b0000000110000000, 16'b1111011110100100, 16'b1111111111111111, 16'b1111111101100101, 16'b1111111000100011, 16'b1111111111101100, 16'b0000000000000000, 16'b0000010001100001, 16'b1111111110100110, 16'b1111111111010011, 16'b0000000010101000, 16'b1111101010110110, 16'b0000000000110001, 16'b1111110001111110, 16'b0000010111000111, 16'b1111111110010100, 16'b1111111000110000, 16'b1111101110011111, 16'b1111111111101010, 16'b1111101001010110, 16'b1111100110000101, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000111110011, 16'b1111111111100011, 16'b1111110110011101, 16'b1111111101101011, 16'b1111111111010000, 16'b0000000000000000, 16'b1111111110111111, 16'b1111101001100110}
};

localparam logic signed [15:0] bias [32] = '{
16'b0000001000011100,  // 0.5280959606170654
16'b0000001101011101,  // 0.8414360880851746
16'b0000000110010111,  // 0.397830605506897
16'b0000000110100100,  // 0.4105983078479767
16'b1111000101011110,  // -3.657735586166382
16'b1111110001101000,  // -0.8977976441383362
16'b0000011011010010,  // 1.7051936388015747
16'b1111101011100100,  // -1.2765135765075684
16'b1111110110101010,  // -0.5837795734405518
16'b0000101011001100,  // 2.699671983718872
16'b0000000011011110,  // 0.2170683741569519
16'b0000001110000110,  // 0.8814588785171509
16'b1111010101110110,  // -2.634300947189331
16'b1111100001111101,  // -1.877297282218933
16'b0000011010100110,  // 1.6625694036483765
16'b0000101011111011,  // 2.7459704875946045
16'b1111111000010110,  // -0.47838035225868225
16'b0000011011001011,  // 1.6984987258911133
16'b0000001101101011,  // 0.8548859357833862
16'b0000010000000100,  // 1.0045719146728516
16'b0000010110101101,  // 1.4197649955749512
16'b0000001101010100,  // 0.832463800907135
16'b0000001000101100,  // 0.5434179306030273
16'b0000001110110101,  // 0.9277304410934448
16'b1111111010100001,  // -0.3426123857498169
16'b1111110111000011,  // -0.5587119460105896
16'b1111110110000100,  // -0.6208624839782715
16'b1111101011100001,  // -1.2802538871765137
16'b0000000000111100,  // 0.05940237268805504
16'b1111110010110110,  // -0.8213341236114502
16'b0000001110000011,  // 0.8783953189849854
16'b1111110000110011   // -0.949700653553009
};
endpackage