// Width: 14
// NFRAC: 7
package dense_3_14_7;

localparam logic signed [13:0] weights [32][32] = '{ 
{14'b11111111111001, 14'b11111111001000, 14'b11111111001100, 14'b11111111100111, 14'b00000000101011, 14'b00000000000101, 14'b11111111111110, 14'b11111111111111, 14'b11111111111111, 14'b11111111111111, 14'b00000000010000, 14'b11111110111100, 14'b11111111111000, 14'b00000001101100, 14'b11111111100001, 14'b11111110001000, 14'b11111111111011, 14'b00000000001110, 14'b00000000110111, 14'b11111111010011, 14'b11111101110111, 14'b11111111111010, 14'b00000000000110, 14'b11111111001100, 14'b00000000000000, 14'b00000010000001, 14'b11111101000101, 14'b11111111100011, 14'b11111111001110, 14'b11111111101100, 14'b00000000110110, 14'b11111111101011}, 
{14'b00000001011111, 14'b00000011011101, 14'b00000000110011, 14'b11111110101011, 14'b00000000011111, 14'b11111111011101, 14'b11111111110010, 14'b00000010001011, 14'b00000000000000, 14'b11111111111111, 14'b11111111111011, 14'b11111110110100, 14'b11111111100110, 14'b00000001000101, 14'b11111011110010, 14'b11111111000011, 14'b11111111111111, 14'b11111111111110, 14'b11111111111001, 14'b11111111101010, 14'b11111111011110, 14'b11111111011100, 14'b00000000000010, 14'b11111111111111, 14'b11111111111111, 14'b11111101110110, 14'b00000000000001, 14'b00000000111100, 14'b11111111110111, 14'b11111110100111, 14'b00000000000000, 14'b00000000000100}, 
{14'b11111110000001, 14'b00000000010111, 14'b00000000000001, 14'b00000000101001, 14'b11111110101111, 14'b00000000000000, 14'b00000000000000, 14'b11111110010100, 14'b00000001000100, 14'b11111111011110, 14'b11111111011110, 14'b11111101000001, 14'b11111111011000, 14'b00000001000001, 14'b00000000100001, 14'b11111111111111, 14'b11111111110001, 14'b11111111111100, 14'b11111110010111, 14'b00000000000000, 14'b00000000001111, 14'b00000000001000, 14'b00000000011010, 14'b00000001110000, 14'b00000000000100, 14'b11111110011011, 14'b00000001100010, 14'b00000000000000, 14'b00000000010101, 14'b11111111111101, 14'b00000000000000, 14'b00000100100010}, 
{14'b00000001101011, 14'b11111111111111, 14'b11111111100111, 14'b00000010100111, 14'b00000010011101, 14'b00000000000000, 14'b00000000001001, 14'b00000001101000, 14'b11111111001101, 14'b11111111111111, 14'b11111110010110, 14'b00000000001111, 14'b00000000100010, 14'b11111110100000, 14'b00000000001011, 14'b11111111101011, 14'b11111111111111, 14'b11111111010001, 14'b00000000000100, 14'b00000000000111, 14'b00000000000010, 14'b11111111110110, 14'b00000010011000, 14'b00000001010111, 14'b00000001010100, 14'b00000000111111, 14'b00000001010111, 14'b00000000000000, 14'b11111111110000, 14'b00000001110011, 14'b00000000111111, 14'b11111111101001}, 
{14'b00000010000000, 14'b11111111110100, 14'b11111110100111, 14'b11111100111111, 14'b00000001111010, 14'b00000000000000, 14'b11111110010110, 14'b11111110110111, 14'b11111111110100, 14'b11111100110000, 14'b11111011100101, 14'b00000001111001, 14'b00000010101011, 14'b00000010000101, 14'b11111101101100, 14'b11111100111001, 14'b00000000000000, 14'b11111111011011, 14'b00000000110011, 14'b00000000100011, 14'b11111111001111, 14'b11111111111110, 14'b00000010111000, 14'b11111010100000, 14'b00000000010110, 14'b11111101010111, 14'b00000000010000, 14'b11111111000000, 14'b11111110110011, 14'b11111111111111, 14'b00000000010001, 14'b00000010010100}, 
{14'b00000000001011, 14'b11111111110101, 14'b11111110110001, 14'b11111110111101, 14'b00000001011111, 14'b00000000000000, 14'b11111110111000, 14'b11111111011101, 14'b11111110010010, 14'b11111111101111, 14'b11111111111111, 14'b00000000101001, 14'b00000000000000, 14'b00000001011011, 14'b11111101111110, 14'b11111111011111, 14'b00000000010110, 14'b11111110110100, 14'b11111111001101, 14'b11111111111111, 14'b00000000000011, 14'b00000001001100, 14'b00000001110111, 14'b11111111111101, 14'b11111111111111, 14'b00000001100110, 14'b11111101110011, 14'b11111111111111, 14'b11111111000011, 14'b11111111110110, 14'b11111111111111, 14'b00000000000001}, 
{14'b00000000010000, 14'b11111110101010, 14'b00000000011011, 14'b11111111110110, 14'b11111111111110, 14'b00000000100110, 14'b11111111100100, 14'b11111101010010, 14'b11111111111111, 14'b11111111001010, 14'b11111110001011, 14'b00000001111000, 14'b00000000000001, 14'b00000010101111, 14'b00000011010100, 14'b00000000000000, 14'b11111111111111, 14'b11111110101111, 14'b11111111110000, 14'b00000001000101, 14'b11111100111111, 14'b00000000100111, 14'b00000001010011, 14'b00000000000100, 14'b00000000100110, 14'b00000100111110, 14'b11111110011011, 14'b11111111101000, 14'b11111111001111, 14'b00000001111100, 14'b11111111110011, 14'b11111111010100}, 
{14'b11111101100111, 14'b00000000000110, 14'b11111101011110, 14'b00000001101111, 14'b00000100000111, 14'b00000000011101, 14'b00000000000000, 14'b00000000001100, 14'b11111111111111, 14'b00000000100000, 14'b00000101001101, 14'b11111111111111, 14'b00000001100001, 14'b00000010011111, 14'b00000011000100, 14'b00000100001100, 14'b00000000000000, 14'b11111110000101, 14'b00000001010110, 14'b11111111111110, 14'b11111101011100, 14'b11111111000101, 14'b00000000000011, 14'b11111111101010, 14'b11111101111111, 14'b00000111100000, 14'b11111111000111, 14'b00000000000000, 14'b00000000000000, 14'b00000011100010, 14'b00000000010110, 14'b00000001100100}, 
{14'b00000001101100, 14'b11111111111011, 14'b00000000000000, 14'b11111111110100, 14'b00000000010100, 14'b11111111110110, 14'b11111111111111, 14'b00000000101000, 14'b00000000110110, 14'b11111110111001, 14'b00000000100011, 14'b00000000101111, 14'b00000000000011, 14'b00000001010101, 14'b11111111000110, 14'b11111100110011, 14'b00000000000000, 14'b11111111111100, 14'b11111111111001, 14'b11111110000000, 14'b11111111111111, 14'b00000000000000, 14'b11111111001100, 14'b11111111111100, 14'b11111111100111, 14'b00000000100111, 14'b00000001011111, 14'b11111111100001, 14'b11111111110011, 14'b11111111110101, 14'b00000000000110, 14'b11111110011011}, 
{14'b11111111010010, 14'b00000001100010, 14'b00000000000000, 14'b00000000000000, 14'b00000011001010, 14'b00000001010010, 14'b11111111111111, 14'b11111101110001, 14'b00000000011110, 14'b11111101001101, 14'b11111010011000, 14'b11111111111111, 14'b00000000000000, 14'b00000001101101, 14'b00000000011100, 14'b00000000000000, 14'b11111110101011, 14'b00000000000000, 14'b00000000000001, 14'b00000000001111, 14'b00000000111110, 14'b11111111111001, 14'b11111110100011, 14'b00000000000010, 14'b11111111111101, 14'b00000100010100, 14'b00000001010011, 14'b11111111111111, 14'b11111111101101, 14'b00000010101011, 14'b11111111110101, 14'b11111111101001}, 
{14'b11111101111010, 14'b00000000101100, 14'b11111111110111, 14'b11111111111111, 14'b11111111000000, 14'b11111110011111, 14'b00000000001100, 14'b00000000100100, 14'b11111111111111, 14'b11111111010100, 14'b11111101101101, 14'b00000000110011, 14'b00000001001101, 14'b00000000000000, 14'b00000011010110, 14'b11111101110000, 14'b00000000011010, 14'b11111110011011, 14'b00000001001000, 14'b11111111111111, 14'b11111111110110, 14'b00000000010001, 14'b00000000011111, 14'b00000000000000, 14'b11111110000001, 14'b00000000000111, 14'b11111101110000, 14'b11111111110101, 14'b11111111111111, 14'b00000010101100, 14'b11111111001111, 14'b00000000000000}, 
{14'b11111111111111, 14'b00000000011101, 14'b00000000000000, 14'b00000001100100, 14'b11111111100010, 14'b11111111110100, 14'b00000000001110, 14'b11111111111110, 14'b11111111110100, 14'b00000010100100, 14'b00000010110010, 14'b00000000000000, 14'b11111110101010, 14'b11111101001100, 14'b11111111110011, 14'b00000000000000, 14'b00000000000000, 14'b11111111101111, 14'b11111110000110, 14'b00000001100001, 14'b00000000000000, 14'b00000001011110, 14'b11111111111111, 14'b00000010001111, 14'b00000000011111, 14'b00000001001110, 14'b00000001110100, 14'b11111111110010, 14'b11111110011011, 14'b11111110001111, 14'b11111111111110, 14'b11111101010100}, 
{14'b11111111000110, 14'b11111111111111, 14'b00000000011110, 14'b11111110010100, 14'b00000000010110, 14'b11111111111111, 14'b11111111001000, 14'b11111111111101, 14'b11111111011111, 14'b00000000001001, 14'b00000000010011, 14'b11111111101101, 14'b00000000000100, 14'b00000000110000, 14'b11111101011111, 14'b11111111000001, 14'b00000000111010, 14'b11111111010010, 14'b00000000000000, 14'b11111111111001, 14'b00000000110001, 14'b00000000000010, 14'b11111111111000, 14'b00000000001010, 14'b00000001000100, 14'b11111111100101, 14'b00000000000000, 14'b11111110001100, 14'b11111111001101, 14'b11111111111110, 14'b00000000101100, 14'b00000000000000}, 
{14'b11111101111010, 14'b00000001101011, 14'b11111111111111, 14'b11111111111110, 14'b11111111111101, 14'b00000000101100, 14'b11111111111111, 14'b00000011000101, 14'b11111111111100, 14'b11111111111111, 14'b00000000110100, 14'b00000000001010, 14'b00000000000001, 14'b00000000000000, 14'b00000000011111, 14'b00000001010100, 14'b00000000101101, 14'b00000000101010, 14'b11111111111101, 14'b00000001001110, 14'b00000000011001, 14'b00000000001010, 14'b11111111111101, 14'b00000001000001, 14'b11111111100110, 14'b11111110101001, 14'b11111111101000, 14'b11111111111111, 14'b00000000011010, 14'b00000000000111, 14'b00000000110010, 14'b00000001111010}, 
{14'b11111111111011, 14'b11111110011100, 14'b00000000001101, 14'b11111111111111, 14'b00000011101010, 14'b11111111001010, 14'b11111101101101, 14'b00000000000000, 14'b00000000000000, 14'b11111111111001, 14'b00000000001100, 14'b00000001101111, 14'b00000001010010, 14'b00000000000010, 14'b00000000001000, 14'b11111111010011, 14'b00000000001000, 14'b11111111110110, 14'b00000000000000, 14'b00000000010011, 14'b11111111110110, 14'b00000000000100, 14'b00000001000100, 14'b00000000001001, 14'b11111111111100, 14'b11111110010110, 14'b00000000110100, 14'b11111111111111, 14'b11111111111111, 14'b11111111100100, 14'b11111111111010, 14'b11111111101111}, 
{14'b00000000000001, 14'b11111111101111, 14'b11111111011111, 14'b11111111001000, 14'b11111101110100, 14'b00000010011100, 14'b00000000000000, 14'b00000000101011, 14'b00000001001001, 14'b00000000000011, 14'b11111111110111, 14'b00000001111001, 14'b00000000111001, 14'b11111110100010, 14'b11111111010110, 14'b11111111110101, 14'b11111110011010, 14'b11111111111011, 14'b00000000000000, 14'b11111111111110, 14'b00000000100111, 14'b11111111011100, 14'b00000000000000, 14'b00000000010011, 14'b11111111111111, 14'b11111110101000, 14'b00000000101000, 14'b00000000000000, 14'b00000000001011, 14'b00000000000010, 14'b11111110101111, 14'b00000000000101}, 
{14'b11111111001101, 14'b11111111010111, 14'b00000000010011, 14'b11111111100000, 14'b11111111101001, 14'b00000000011101, 14'b11111111111110, 14'b00000000001000, 14'b00000000100001, 14'b11111111111111, 14'b00000000011111, 14'b11111111011111, 14'b11111111111101, 14'b11111111111111, 14'b00000000011010, 14'b11111111111111, 14'b00000001111101, 14'b11111111111011, 14'b00000000111111, 14'b11111111010100, 14'b00000000101000, 14'b00000000010000, 14'b00000000010101, 14'b00000000001001, 14'b11111111101011, 14'b11111110111000, 14'b11111110111101, 14'b00000000011011, 14'b11111111101010, 14'b00000000000000, 14'b11111111111000, 14'b00000000111011}, 
{14'b11111111111111, 14'b11111110011000, 14'b11111110011010, 14'b11111111111111, 14'b00000010100001, 14'b11111111101000, 14'b00000000000000, 14'b00000001111011, 14'b11111111011010, 14'b00000000000000, 14'b11111110010101, 14'b11111110000010, 14'b00000001110010, 14'b00000000100110, 14'b11111111100000, 14'b11111110111001, 14'b00000000101100, 14'b00000000000000, 14'b11111111000011, 14'b00000000000110, 14'b00000000010001, 14'b11111111101001, 14'b00000001001000, 14'b11111100000101, 14'b00000000001010, 14'b00000000111101, 14'b11111111110101, 14'b00000000000011, 14'b11111111000100, 14'b11111111111111, 14'b11111111001100, 14'b11111111111001}, 
{14'b00000000110110, 14'b00000001011000, 14'b00000010001100, 14'b11111111001011, 14'b00000001101010, 14'b00000001001110, 14'b00000000000000, 14'b00000001110100, 14'b00000001011011, 14'b11111111100100, 14'b00000010110011, 14'b11111110100110, 14'b00000010011111, 14'b00000001110010, 14'b11111011101101, 14'b11111111111111, 14'b00000000000000, 14'b00000000000001, 14'b00000001000010, 14'b11111101111111, 14'b00000000111000, 14'b11111111001001, 14'b11111110000010, 14'b11111111010111, 14'b00000001010100, 14'b11111101010111, 14'b11111110101011, 14'b11111111110101, 14'b11111111111111, 14'b11111101101111, 14'b00000001100101, 14'b00000000000000}, 
{14'b11111111110011, 14'b00000000000000, 14'b11111111111111, 14'b11111111111111, 14'b11111110100110, 14'b00000000000010, 14'b00000000000010, 14'b11111111111100, 14'b11111111111001, 14'b11111111110100, 14'b00000000100011, 14'b11111111111111, 14'b00000000010101, 14'b11111110101000, 14'b00000000011011, 14'b11111111111111, 14'b00000000100100, 14'b00000001110010, 14'b11111110100101, 14'b00000000001101, 14'b11111111100110, 14'b00000000100000, 14'b00000000110000, 14'b11111111101010, 14'b11111110111111, 14'b00000000000101, 14'b00000011010100, 14'b11111111111001, 14'b11111111111100, 14'b00000001010011, 14'b00000000000000, 14'b00000011011100}, 
{14'b11111101111010, 14'b00000000001001, 14'b11111111001000, 14'b00000001100010, 14'b00000000011100, 14'b11111111110111, 14'b11111111111111, 14'b11111111111111, 14'b11111110110010, 14'b11111111110111, 14'b00000000000000, 14'b11111101110001, 14'b00000000000011, 14'b11111111110101, 14'b11111111111111, 14'b11111111111111, 14'b11111111100010, 14'b00000000000001, 14'b00000000000000, 14'b00000000101000, 14'b00000000000100, 14'b00000000000000, 14'b00000000000000, 14'b11111111111101, 14'b00000000000000, 14'b00000000000100, 14'b00000010010100, 14'b11111111111111, 14'b11111111111111, 14'b11111111110101, 14'b00000000101100, 14'b11111111111001}, 
{14'b11111111111111, 14'b11111111011001, 14'b00000000110100, 14'b00000000001010, 14'b11111110100000, 14'b00000000000000, 14'b00000001001001, 14'b11111111111111, 14'b00000000000000, 14'b11111111100110, 14'b00000000011101, 14'b00000000000100, 14'b00000001010010, 14'b11111101110011, 14'b11111111100111, 14'b11111111111011, 14'b00000000110111, 14'b11111110011101, 14'b00000000000101, 14'b11111100111110, 14'b11111111111011, 14'b11111111100001, 14'b11111111110101, 14'b00000001001011, 14'b11111111101100, 14'b11111110111000, 14'b00000000010111, 14'b00000000000000, 14'b00000001100101, 14'b00000010000101, 14'b11111110101100, 14'b11111110001101}, 
{14'b00000000010001, 14'b00000000000110, 14'b11111110010101, 14'b11111111110001, 14'b11111111111111, 14'b00000000000000, 14'b00000000011011, 14'b00000001101001, 14'b00000000000000, 14'b00000000000101, 14'b00000000010001, 14'b11111101110101, 14'b11111111101110, 14'b11111101100101, 14'b00000001111011, 14'b00000000000000, 14'b11111111111111, 14'b11111101011011, 14'b11111111111111, 14'b11111111101100, 14'b11111111111010, 14'b00000000000000, 14'b00000000001111, 14'b11111111011001, 14'b00000000001101, 14'b00000001101001, 14'b00000001101101, 14'b00000001100011, 14'b00000001001110, 14'b00000000000000, 14'b00000000011101, 14'b00000011001000}, 
{14'b11111111111001, 14'b11111111000011, 14'b00000001100011, 14'b11111111100101, 14'b00000000010001, 14'b00000000101010, 14'b11111111111111, 14'b11111110110110, 14'b11111111101010, 14'b11111101100110, 14'b00000001110010, 14'b00000000000000, 14'b00000001101011, 14'b00000010101011, 14'b11111111100010, 14'b11111100100001, 14'b11111111100101, 14'b00000001111000, 14'b11111110110111, 14'b11111111001010, 14'b00000000001111, 14'b00000000000000, 14'b11111101110100, 14'b11111111001111, 14'b11111111110101, 14'b11111111100000, 14'b00000000011100, 14'b00000010110100, 14'b00000000111110, 14'b11111111111111, 14'b00000000010100, 14'b00000000000111}, 
{14'b00000000001010, 14'b00000001110100, 14'b00000000000000, 14'b00000001001011, 14'b00000011010100, 14'b11111111010100, 14'b11111111111111, 14'b11111111110100, 14'b00000001001011, 14'b11111111001110, 14'b11111111111111, 14'b00000001010101, 14'b00000000000010, 14'b00000000000111, 14'b11111001111001, 14'b11111111101011, 14'b00000000000000, 14'b00000000110011, 14'b11111111111111, 14'b00000001001100, 14'b11111111111111, 14'b11111111010011, 14'b11111101110000, 14'b00000000100001, 14'b00000001001001, 14'b11111011100100, 14'b11111111111111, 14'b00000000000000, 14'b00000010001011, 14'b11111100110010, 14'b00000000000000, 14'b11111111111110}, 
{14'b00000000000010, 14'b11111110101001, 14'b00000000001101, 14'b11111111111100, 14'b00000000001101, 14'b00000010000111, 14'b11111101000110, 14'b00000000001000, 14'b00000001101100, 14'b11111110101001, 14'b11111111111010, 14'b00000000001100, 14'b11111111111101, 14'b00000000101101, 14'b00000000011011, 14'b11111111111011, 14'b00000000010001, 14'b00000000000000, 14'b00000000000101, 14'b00000001100001, 14'b11111111111000, 14'b11111110000100, 14'b11111101100101, 14'b11111111001110, 14'b11111101101000, 14'b00000000110101, 14'b00000010011111, 14'b00000001011110, 14'b11111111111101, 14'b11111110100000, 14'b11111110110000, 14'b00000000001111}, 
{14'b00000000001101, 14'b11111110000101, 14'b11111111111011, 14'b00000000100110, 14'b11111110000101, 14'b00000000101011, 14'b11111111111111, 14'b11111111111111, 14'b11111111111111, 14'b00000000000000, 14'b00000001000011, 14'b11111111111011, 14'b00000000000010, 14'b00000000000000, 14'b00000000100000, 14'b11111111111011, 14'b00000000000000, 14'b11111111111111, 14'b11111110101101, 14'b11111101111110, 14'b11111111111111, 14'b11111101110111, 14'b11111110110010, 14'b11111110100000, 14'b00000011100011, 14'b00000000000100, 14'b11111111110100, 14'b00000001010001, 14'b00000011100101, 14'b00000001100101, 14'b11111011110000, 14'b11111111010000}, 
{14'b00000001100000, 14'b11111111111111, 14'b00000001000000, 14'b11111111111010, 14'b00000001111011, 14'b11111111011011, 14'b00000000010010, 14'b00000001101011, 14'b00000001000100, 14'b11111101111010, 14'b11111111110000, 14'b00000000011111, 14'b00000000010001, 14'b11111111111100, 14'b00000000010101, 14'b00000000000000, 14'b00000001011100, 14'b00000000001000, 14'b00000001011111, 14'b11111111101111, 14'b11111111011111, 14'b11111111101100, 14'b11111111111111, 14'b00000001001101, 14'b11111111001100, 14'b11111111111110, 14'b00000000000000, 14'b00000000000000, 14'b00000000000000, 14'b00000001001010, 14'b11111110101101, 14'b11111111111010}, 
{14'b11111111111111, 14'b11111111111000, 14'b11111110001000, 14'b00000001001000, 14'b00000000111001, 14'b11111111100011, 14'b11111111111111, 14'b11111111000101, 14'b00000000000001, 14'b11111111111111, 14'b11111110110010, 14'b11111111000000, 14'b00000001111010, 14'b00000000000000, 14'b11111111011111, 14'b11111111111111, 14'b00000000110110, 14'b11111111111111, 14'b11111111111111, 14'b11111111001000, 14'b00000001010000, 14'b00000000000000, 14'b00000000100111, 14'b11111111111000, 14'b00000000101000, 14'b00000000000000, 14'b00000000000000, 14'b00000000111101, 14'b11111111001110, 14'b11111111110100, 14'b00000000101001, 14'b11111111100100}, 
{14'b11111111111011, 14'b11111110110001, 14'b00000010011000, 14'b11111111101111, 14'b00000000110010, 14'b11111110110110, 14'b00000000000000, 14'b00000000001000, 14'b11111110000101, 14'b11111111111100, 14'b11111111100000, 14'b00000000001110, 14'b11111110101100, 14'b00000000100011, 14'b00000000110011, 14'b00000000011100, 14'b00000000010101, 14'b11111111110110, 14'b11111101001010, 14'b11111111111100, 14'b11111111110001, 14'b00000000100011, 14'b11111111100011, 14'b11111111111111, 14'b00000000110010, 14'b11111111110100, 14'b11111111111100, 14'b00000001100011, 14'b11111110011010, 14'b11111110110100, 14'b00000001011001, 14'b00000000001001}, 
{14'b00000001101110, 14'b00000000110011, 14'b00000000000000, 14'b11111111010111, 14'b11111111101011, 14'b11111111111111, 14'b00000000000000, 14'b11111111101110, 14'b11111111100000, 14'b11111111100001, 14'b00000000000000, 14'b00000000101000, 14'b00000000000001, 14'b00000000001101, 14'b11111111110100, 14'b00000000000001, 14'b11111111011000, 14'b00000000000000, 14'b11111111111011, 14'b11111111111111, 14'b00000000000000, 14'b00000000001111, 14'b00000000011000, 14'b00000000000000, 14'b00000000000000, 14'b11111101100011, 14'b11111111001100, 14'b00000000000001, 14'b00000000000101, 14'b00000000000000, 14'b11111111010010, 14'b00000000000101}, 
{14'b00000000110000, 14'b11111011110100, 14'b11111111111111, 14'b11111111101100, 14'b11111111000100, 14'b11111111111101, 14'b00000000000000, 14'b00000010001100, 14'b11111111110100, 14'b11111111111010, 14'b00000000010101, 14'b11111101010110, 14'b00000000000110, 14'b11111110001111, 14'b00000010111000, 14'b11111111110010, 14'b11111111000110, 14'b11111101110011, 14'b11111111111101, 14'b11111101001010, 14'b11111100110000, 14'b11111111111111, 14'b00000000000000, 14'b00000000000000, 14'b00000000111110, 14'b11111111111100, 14'b11111110110011, 14'b11111111101101, 14'b11111111111010, 14'b00000000000000, 14'b11111111110111, 14'b11111101001100}
};

localparam logic signed [13:0] bias [32] = '{
14'b00000001000011,  // 0.5280959606170654
14'b00000001101011,  // 0.8414360880851746
14'b00000000110010,  // 0.397830605506897
14'b00000000110100,  // 0.4105983078479767
14'b11111000101011,  // -3.657735586166382
14'b11111110001101,  // -0.8977976441383362
14'b00000011011010,  // 1.7051936388015747
14'b11111101011100,  // -1.2765135765075684
14'b11111110110101,  // -0.5837795734405518
14'b00000101011001,  // 2.699671983718872
14'b00000000011011,  // 0.2170683741569519
14'b00000001110000,  // 0.8814588785171509
14'b11111010101110,  // -2.634300947189331
14'b11111100001111,  // -1.877297282218933
14'b00000011010100,  // 1.6625694036483765
14'b00000101011111,  // 2.7459704875946045
14'b11111111000010,  // -0.47838035225868225
14'b00000011011001,  // 1.6984987258911133
14'b00000001101101,  // 0.8548859357833862
14'b00000010000000,  // 1.0045719146728516
14'b00000010110101,  // 1.4197649955749512
14'b00000001101010,  // 0.832463800907135
14'b00000001000101,  // 0.5434179306030273
14'b00000001110110,  // 0.9277304410934448
14'b11111111010100,  // -0.3426123857498169
14'b11111110111000,  // -0.5587119460105896
14'b11111110110000,  // -0.6208624839782715
14'b11111101011100,  // -1.2802538871765137
14'b00000000000111,  // 0.05940237268805504
14'b11111110010110,  // -0.8213341236114502
14'b00000001110000,  // 0.8783953189849854
14'b11111110000110   // -0.949700653553009
};
endpackage