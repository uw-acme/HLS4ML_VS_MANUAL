// Width: 11
// NFRAC: 5
package dense_4_11_5;

localparam logic signed [10:0] weights [32][5] = '{ 
{11'b11111111111, 11'b00000001010, 11'b11111110110, 11'b00000000010, 11'b11111111100}, 
{11'b11111101110, 11'b11111111110, 11'b00000001110, 11'b11111111111, 11'b00000000000}, 
{11'b00000001011, 11'b00000000110, 11'b11111111111, 11'b11111110011, 11'b11111111001}, 
{11'b11111110011, 11'b11111110100, 11'b11111111100, 11'b00000001001, 11'b00000000111}, 
{11'b00000000011, 11'b00000000100, 11'b00000000101, 11'b11111111111, 11'b11111011111}, 
{11'b00000001010, 11'b11111110011, 11'b00000000101, 11'b11111111010, 11'b11111111010}, 
{11'b11111110011, 11'b00000000001, 11'b11111111111, 11'b00000000101, 11'b00000000010}, 
{11'b11111111111, 11'b00000001001, 11'b11111110011, 11'b00000000101, 11'b00000000100}, 
{11'b00000000101, 11'b11111111010, 11'b00000000000, 11'b11111110001, 11'b11111111000}, 
{11'b11111111111, 11'b11111110111, 11'b00000000101, 11'b00000001101, 11'b00000000000}, 
{11'b11111111011, 11'b11111111011, 11'b00000000000, 11'b00000010010, 11'b11111110111}, 
{11'b00000000101, 11'b00000000111, 11'b11111110101, 11'b11111111111, 11'b00000000011}, 
{11'b00000000000, 11'b00000000101, 11'b00000000000, 11'b11111111001, 11'b11111101100}, 
{11'b00000000101, 11'b00000000010, 11'b00000001101, 11'b11111111101, 11'b11111110010}, 
{11'b00000000010, 11'b11111111110, 11'b11111110100, 11'b11111111110, 11'b00000010001}, 
{11'b11111110000, 11'b11111111000, 11'b11111111000, 11'b00000001100, 11'b00000000001}, 
{11'b00000001011, 11'b11111111010, 11'b11111111011, 11'b11111111000, 11'b11111111110}, 
{11'b00000000110, 11'b11111111110, 11'b11111110010, 11'b11111111111, 11'b00000000010}, 
{11'b00000001000, 11'b00000000001, 11'b11111111001, 11'b00000000000, 11'b11111110011}, 
{11'b00000000111, 11'b11111111101, 11'b11111111001, 11'b00000000110, 11'b00000000011}, 
{11'b00000000010, 11'b11111111111, 11'b00000001001, 11'b11111110010, 11'b11111111111}, 
{11'b00000000000, 11'b00000000011, 11'b00000001111, 11'b11111101111, 11'b11111101100}, 
{11'b11111111100, 11'b00000000011, 11'b00000000101, 11'b11111110100, 11'b00000010000}, 
{11'b11111111111, 11'b00000000101, 11'b00000001001, 11'b00000000001, 11'b11111101101}, 
{11'b11111111010, 11'b00000001011, 11'b11111111000, 11'b00000000000, 11'b00000001100}, 
{11'b00000000000, 11'b00000001000, 11'b00000000000, 11'b11111101000, 11'b00000010001}, 
{11'b11111110001, 11'b11111111000, 11'b00000000110, 11'b00000000111, 11'b00000000110}, 
{11'b00000000000, 11'b00000000111, 11'b11111111110, 11'b11111111011, 11'b00000000001}, 
{11'b11111111100, 11'b00000000111, 11'b11111101111, 11'b00000000100, 11'b11111111010}, 
{11'b11111111111, 11'b00000000100, 11'b11111111010, 11'b11111110011, 11'b00000010010}, 
{11'b00000001110, 11'b00000000010, 11'b00000001010, 11'b11111101101, 11'b11111110101}, 
{11'b11111111110, 11'b11111110011, 11'b00000001011, 11'b00000000010, 11'b00000000100}
};

localparam logic signed [10:0] bias [5] = '{
11'b11111111110,  // -0.06223141402006149
11'b11111111101,  // -0.06270556896924973
11'b11111111101,  // -0.07014333456754684
11'b00000000010,  // 0.0820775106549263
11'b00000000110   // 0.2155742198228836
};
endpackage