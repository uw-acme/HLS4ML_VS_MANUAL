// Width: 22
// NFRAC: 11
package dense_1_22_11;

localparam logic signed [21:0] weights [16][64] = '{ 
{22'b0000000000001000001010, 22'b1111111111101011001001, 22'b1111111111111010001101, 22'b1111111111111000110000, 22'b1111111111110011000010, 22'b0000000000000011100010, 22'b1111111111011110110100, 22'b0000000000000000000000, 22'b0000000000000001110110, 22'b0000000000001000011011, 22'b0000000000000000000110, 22'b1111111111110011000011, 22'b1111111111111111111101, 22'b0000000000000110101100, 22'b0000000000000001000100, 22'b1111111111110111101000, 22'b0000000000000111011100, 22'b0000000000000001111000, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b0000000000001100000011, 22'b1111111111110101011001, 22'b1111111111111111010010, 22'b0000000000001111001000, 22'b1111111111110101101101, 22'b1111111111101010001010, 22'b1111111111110111001011, 22'b1111111111111001110000, 22'b1111111111111100101001, 22'b1111111111111111111100, 22'b0000000000000001001101, 22'b0000000000000111110110, 22'b0000000000000110010000, 22'b1111111111111111100101, 22'b0000000000000000000000, 22'b0000000000001001111101, 22'b1111111111111111011011, 22'b1111111111110111111101, 22'b0000000000000000110111, 22'b0000000000000110001010, 22'b1111111111111111100111, 22'b0000000000001000110011, 22'b1111111111110111011110, 22'b0000000000011101101110, 22'b1111111111111111111101, 22'b0000000000001110011110, 22'b0000000000000000000000, 22'b0000000000000101111001, 22'b0000000000000110010001, 22'b1111111111111111001111, 22'b0000000000000000000000, 22'b0000000000000101001000, 22'b0000000000000110111010, 22'b0000000000000010011111, 22'b1111111111111100010011, 22'b1111111111110110000100, 22'b0000000000010001001010, 22'b1111111111110000000000, 22'b0000000000001110111101, 22'b1111111111110100101010, 22'b0000000000011001011000, 22'b1111111111111111110000, 22'b0000000000000000010111, 22'b0000000000000010100110}, 
{22'b0000000000000000000101, 22'b1111111111110101101111, 22'b1111111111111011110000, 22'b1111111111110111000011, 22'b1111111111110101110101, 22'b0000000000000011011010, 22'b1111111111100111110110, 22'b1111111111111111111011, 22'b1111111111111000101110, 22'b0000000000000101100001, 22'b0000000000000000001101, 22'b1111111111111101001111, 22'b0000000000000110010011, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b0000000000000110101001, 22'b1111111111111111110011, 22'b0000000000000000000000, 22'b1111111111111010001010, 22'b1111111111110111111111, 22'b0000000000001110001001, 22'b1111111111111101011010, 22'b0000000000000001100010, 22'b0000000000010110010111, 22'b0000000000001000001111, 22'b1111111111111000101000, 22'b1111111111111000100111, 22'b1111111111111111111111, 22'b1111111111111100110000, 22'b1111111111110011000001, 22'b1111111111111110000101, 22'b0000000000001110100011, 22'b0000000000001000111010, 22'b0000000000010001100110, 22'b0000000000010100001000, 22'b0000000000000001100111, 22'b1111111111111100001101, 22'b1111111111110010000111, 22'b0000000000000001110100, 22'b0000000000000110000010, 22'b0000000000000000101110, 22'b0000000000000110100110, 22'b1111111111111001001100, 22'b0000000000001000000100, 22'b0000000000000101100000, 22'b0000000000000001100110, 22'b1111111111110101000111, 22'b0000000000000010100010, 22'b0000000000001000010101, 22'b0000000000000000111101, 22'b0000000000000000110010, 22'b0000000000100101000010, 22'b1111111111111101100110, 22'b1111111111111100110111, 22'b1111111111111110010000, 22'b1111111111111111110000, 22'b0000000000001000001110, 22'b1111111111110100001010, 22'b0000000000011111100001, 22'b0000000000000000001001, 22'b0000000000010000101010, 22'b0000000000000111101011, 22'b0000000000011010010100, 22'b0000000000000100100000}, 
{22'b1111111111111111110000, 22'b0000000000000000000000, 22'b1111111111111101010101, 22'b1111111111111010010111, 22'b1111111111111010000101, 22'b0000000000000001010101, 22'b0000000000101111011000, 22'b1111111111111111111111, 22'b1111111111010111011111, 22'b1111111111111111111111, 22'b1111111111111111111100, 22'b1111111111111111011011, 22'b1111111111111000101110, 22'b0000000000000000000010, 22'b1111111111111111101100, 22'b0000000000000101011000, 22'b0000000000011100111110, 22'b1111111111111111111111, 22'b0000000000000010010011, 22'b0000000000000000000000, 22'b0000000000001101001100, 22'b1111111111101000111010, 22'b0000000000010010011110, 22'b1111111111101001001010, 22'b0000000000011110010110, 22'b1111111111110100111010, 22'b1111111111111000001010, 22'b1111111111101001000010, 22'b0000000000101000110000, 22'b0000000000001000110100, 22'b0000000000000000010111, 22'b0000000000010000100100, 22'b0000000000100000101001, 22'b1111111111011001110000, 22'b1111111111111100111100, 22'b0000000000000001000001, 22'b1111111111111000100110, 22'b0000000000011100101101, 22'b1111111111111110101111, 22'b0000000000001010000001, 22'b0000000000001010101010, 22'b0000000000001011110101, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b1111111111111111011100, 22'b0000000000000101000001, 22'b1111111111110111000011, 22'b1111111111111010100011, 22'b1111111111111111011100, 22'b0000000000001100100101, 22'b1111111111111010010111, 22'b0000000000000100110011, 22'b1111111111111111111111, 22'b0000000000000100010010, 22'b1111111111111010011000, 22'b1111111111111111111111, 22'b1111111111110110001000, 22'b1111111111101010100100, 22'b1111111111111111111011, 22'b0000000000000000000000, 22'b0000000000110001010111, 22'b0000000000000000011010, 22'b1111111111111111111010, 22'b1111111111110110000110}, 
{22'b1111111111110001010101, 22'b1111111111110100001101, 22'b1111111111101001110101, 22'b0000000000001001110111, 22'b1111111111110101111001, 22'b1111111111010100111010, 22'b1111111111111100010101, 22'b1111111111110110001001, 22'b0000000000000111001010, 22'b1111111111111111111111, 22'b0000000000101000011111, 22'b1111111111111100100111, 22'b1111111111100110111101, 22'b0000000000010010100010, 22'b0000000000000000110011, 22'b1111111111111111111100, 22'b1111111111110001110011, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b1111111111111000110000, 22'b1111111111011011001010, 22'b1111111111111100011011, 22'b1111111111101001101001, 22'b0000000000000110010110, 22'b1111111111110011100111, 22'b1111111111100010100010, 22'b0000000000001010000000, 22'b0000000000010111100100, 22'b0000000000101001011100, 22'b1111111111110001010010, 22'b1111111111101101010110, 22'b0000000000000010010111, 22'b0000000000010000000000, 22'b1111111111100101000101, 22'b1111111111110101111100, 22'b0000000000000000000000, 22'b1111111111101000110001, 22'b0000000000000111110000, 22'b1111111111110001111000, 22'b0000000000000011110100, 22'b0000000000001110101011, 22'b0000000000000101000001, 22'b0000000000000000000000, 22'b0000000000000000101001, 22'b0000000000010001101011, 22'b1111111111111001100110, 22'b1111111111111111111111, 22'b1111111111110100111111, 22'b1111111111111111111111, 22'b1111111111111100111001, 22'b1111111111101100010011, 22'b0000000000000010110001, 22'b1111111111111111111111, 22'b0000000000000110111110, 22'b0000000000001010000101, 22'b0000000000010100101101, 22'b1111111111100001000010, 22'b1111111111100010010001, 22'b1111111111101001011011, 22'b0000000000011011101110, 22'b0000000000110111111110, 22'b1111111111100011001101, 22'b1111111111111110010001, 22'b0000000000001101111001}, 
{22'b0000000000001010111100, 22'b1111111111101100001101, 22'b1111111111110111101100, 22'b1111111111111111111111, 22'b1111111111111011000100, 22'b0000000000001010111000, 22'b0000000000000110000100, 22'b1111111111111111111111, 22'b1111111111101100111000, 22'b1111111111111000010000, 22'b1111111111110100001100, 22'b0000000000000001101100, 22'b0000000000000000000010, 22'b0000000000000000000000, 22'b1111111111111110101101, 22'b0000000000001011011100, 22'b0000000000000100010001, 22'b1111111111110011011011, 22'b0000000000000000111110, 22'b0000000000000000011011, 22'b0000000000000110101110, 22'b1111111111111100001110, 22'b0000000000000010011000, 22'b1111111111111111011000, 22'b0000000000100010000110, 22'b1111111111111010000010, 22'b1111111111110111000000, 22'b1111111111110011000101, 22'b0000000000000000000000, 22'b0000000000000101010001, 22'b0000000000000011101110, 22'b0000000000001000110000, 22'b1111111111111111100110, 22'b0000000000000010010111, 22'b0000000000000100001011, 22'b1111111111111111111111, 22'b0000000000000000001100, 22'b0000000000011100001101, 22'b1111111111110110110000, 22'b1111111111111101100011, 22'b0000000000001101110111, 22'b0000000000000111111101, 22'b1111111111110000010110, 22'b0000000000000000001100, 22'b1111111111011101110100, 22'b1111111111111111111111, 22'b1111111111111100000101, 22'b0000000000000000011000, 22'b1111111111111111111111, 22'b1111111111111111001111, 22'b1111111111111111111111, 22'b0000000000000110000001, 22'b1111111111111111110101, 22'b0000000000001010001010, 22'b1111111111111001111000, 22'b1111111111101000011110, 22'b1111111111110001000100, 22'b1111111111101111101100, 22'b1111111111101100010110, 22'b0000000000010111111001, 22'b0000000000101011111101, 22'b0000000000011001010111, 22'b0000000000000011111011, 22'b1111111111111111111111}, 
{22'b1111111111110001101111, 22'b1111111111101011110100, 22'b0000000000000000000000, 22'b0000000000001001110101, 22'b0000000000001001001000, 22'b1111111111111001001101, 22'b0000000000010010101000, 22'b1111111111111111111111, 22'b0000000000000111110011, 22'b1111111111111111111111, 22'b1111111111111111101100, 22'b1111111111111101101011, 22'b1111111111111010010110, 22'b0000000000010010100000, 22'b1111111111111101001001, 22'b0000000000000000000000, 22'b1111111111101100000000, 22'b1111111111110100101010, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b1111111111111110011110, 22'b1111111111110101111101, 22'b1111111111110101110011, 22'b0000000000001110111001, 22'b1111111111110101110100, 22'b1111111111111111111110, 22'b0000000000001000001100, 22'b1111111111111101101010, 22'b1111111111100010001001, 22'b1111111111111111111111, 22'b1111111111111101110111, 22'b1111111111111111101010, 22'b1111111111111111101000, 22'b0000000000000001010011, 22'b0000000000000100001110, 22'b0000000000001011000100, 22'b0000000000000000011011, 22'b1111111111111100110111, 22'b1111111111110111100110, 22'b1111111111111111111100, 22'b1111111111111010100101, 22'b1111111111101111001111, 22'b0000000000001100110011, 22'b0000000000000000010110, 22'b0000000000010011010011, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b0000000000000011000010, 22'b1111111111110010100101, 22'b0000000000000111011111, 22'b0000000000000000000000, 22'b1111111111111100110001, 22'b1111111111110100011011, 22'b0000000000001100010111, 22'b1111111111111111111111, 22'b0000000000001011000110, 22'b0000000000000110111011, 22'b0000000000000110100001, 22'b1111111111111111011001, 22'b1111111111111111101111, 22'b1111111111100110001000, 22'b1111111111111011111101, 22'b1111111111111110001011, 22'b1111111111111111111111}, 
{22'b1111111111110110111100, 22'b1111111111110101010001, 22'b1111111111110010001100, 22'b1111111111111101110001, 22'b1111111111111011101111, 22'b0000000000000011010101, 22'b1111111111101001101010, 22'b1111111111111011001100, 22'b1111111111111000110100, 22'b1111111111111111111111, 22'b1111111111110110110011, 22'b0000000000001011001000, 22'b0000000000000001001000, 22'b0000000000000100011010, 22'b0000000000001001111110, 22'b0000000000000000000000, 22'b0000000000011001100000, 22'b0000000000000010110111, 22'b0000000000000111110001, 22'b0000000000001000100101, 22'b1111111111111010111111, 22'b0000000000001011101000, 22'b1111111111111000001111, 22'b1111111111101111111100, 22'b0000000000000101100011, 22'b0000000000010000100010, 22'b1111111111111111110111, 22'b0000000000000001101110, 22'b1111111111100001100100, 22'b0000000000001001001010, 22'b0000000000001000100011, 22'b1111111111110100000011, 22'b0000000000001111000101, 22'b0000000000010101010001, 22'b0000000000000000000000, 22'b0000000000001010111101, 22'b1111111111111111111111, 22'b0000000000001001000110, 22'b0000000000000110010111, 22'b0000000000000000000000, 22'b1111111111111100001110, 22'b1111111111110100010111, 22'b0000000000000100100101, 22'b0000000000001111011101, 22'b0000000000010000100111, 22'b1111111111111010100111, 22'b1111111111111101010101, 22'b1111111111111001111011, 22'b1111111111111011101011, 22'b0000000000000011110010, 22'b0000000000000000000110, 22'b0000000000000001000101, 22'b0000000000000000000000, 22'b0000000000000101110011, 22'b1111111111111010011010, 22'b0000000000011000101010, 22'b0000000000001011011001, 22'b1111111111111111001101, 22'b0000000000001100011111, 22'b0000000000000110111100, 22'b1111111111001011111111, 22'b1111111111101101100011, 22'b1111111111111010011111, 22'b1111111111111111101011}, 
{22'b0000000000000000001010, 22'b0000000000000111101001, 22'b1111111111111111111111, 22'b1111111111111111111110, 22'b1111111111110101101100, 22'b1111111111111111000000, 22'b1111111111110111110000, 22'b0000000000000000000000, 22'b0000000000000000111000, 22'b0000000000001100011100, 22'b0000000000000000011101, 22'b1111111111110011111010, 22'b1111111111111101111111, 22'b0000000000000000000000, 22'b1111111111111110010100, 22'b1111111111110001100111, 22'b1111111111100100110110, 22'b1111111111111111111111, 22'b1111111111101100101010, 22'b1111111111110001101110, 22'b1111111111110011100010, 22'b0000000000001011000111, 22'b0000000000000001100000, 22'b1111111111111011011100, 22'b1111111111110010000001, 22'b0000000000000100111110, 22'b0000000000000000000000, 22'b0000000000001111111110, 22'b0000000000011001110010, 22'b1111111111111110101101, 22'b0000000000000000000001, 22'b0000000000000111011000, 22'b1111111111101010001010, 22'b1111111111110100001000, 22'b0000000000000001110001, 22'b0000000000000010111101, 22'b1111111111110111000001, 22'b0000000000000111101010, 22'b0000000000000100001110, 22'b1111111111111011000111, 22'b1111111111110010100100, 22'b1111111111111110110100, 22'b0000000000000001000011, 22'b1111111111111010101011, 22'b0000000000000001110010, 22'b0000000000000111010101, 22'b1111111111111100001011, 22'b0000000000000000110000, 22'b0000000000000000000000, 22'b1111111111111001000001, 22'b1111111111110011100100, 22'b0000000000001101010011, 22'b0000000000000100000011, 22'b1111111111111010010011, 22'b0000000000000100001111, 22'b1111111111111110000001, 22'b1111111111110000110100, 22'b1111111111111011101111, 22'b1111111111111110010101, 22'b1111111111111101110000, 22'b0000000000011010100100, 22'b0000000000000110000110, 22'b1111111111111110011100, 22'b1111111111111111111111}, 
{22'b0000000000000000011110, 22'b0000000000010010110001, 22'b1111111111101101011010, 22'b1111111111111000100110, 22'b0000000000001010010100, 22'b1111111111111001011001, 22'b0000000000100110110000, 22'b1111111111110110110010, 22'b1111111111111111111111, 22'b0000000000001001011000, 22'b0000000000001000001000, 22'b1111111111111111111010, 22'b1111111111111110011101, 22'b1111111111110000100100, 22'b0000000000001001000000, 22'b0000000000000101000111, 22'b1111111111111001110011, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b0000000000001000011111, 22'b1111111111110001010010, 22'b0000000000001100100011, 22'b0000000000010011100111, 22'b1111111111111101001101, 22'b1111111111111111111111, 22'b1111111111111111011110, 22'b1111111111111111111111, 22'b0000000000010111100011, 22'b0000000000000000001010, 22'b1111111111110111010000, 22'b0000000000000000000000, 22'b0000000000001100010010, 22'b1111111111100110000011, 22'b1111111111101110101100, 22'b0000000000000110010111, 22'b0000000000000100011011, 22'b1111111111101101101101, 22'b1111111111111001111100, 22'b1111111111111001001001, 22'b0000000000001100110101, 22'b0000000000001100100000, 22'b0000000000000000000000, 22'b1111111111110111010111, 22'b0000000000000000000001, 22'b0000000000001100101001, 22'b1111111111111110000111, 22'b1111111111111111111111, 22'b0000000000000000010111, 22'b0000000000000111110101, 22'b1111111111111110001010, 22'b1111111111111001110011, 22'b0000000000001011000000, 22'b1111111111111001000111, 22'b0000000000001000111100, 22'b0000000000010010101101, 22'b0000000000000001010001, 22'b0000000000001000011011, 22'b1111111111110011001100, 22'b1111111111110100010000, 22'b0000000000011010100111, 22'b1111111111111011111000, 22'b0000000000000001011110, 22'b1111111111111101000000}, 
{22'b0000000000000000100001, 22'b1111111111110001100001, 22'b0000000000001011110011, 22'b1111111111110110111010, 22'b1111111111111111111001, 22'b0000000000000110110001, 22'b1111111111101101011000, 22'b0000000000000110001000, 22'b0000000000001111101100, 22'b0000000000000100111011, 22'b0000000000001011100110, 22'b0000000000001010010100, 22'b1111111111110110001111, 22'b1111111111111101100100, 22'b1111111111111110010110, 22'b0000000000000000000010, 22'b1111111111100001010010, 22'b0000000000001010010101, 22'b1111111111111110110101, 22'b0000000000000000111111, 22'b1111111111110100101110, 22'b0000000000000010001111, 22'b0000000000000100111001, 22'b1111111111111111111111, 22'b1111111111110001010001, 22'b1111111111111110011110, 22'b1111111111111101011000, 22'b0000000000100111111011, 22'b1111111111101010110011, 22'b0000000000000010001000, 22'b0000000000000011000110, 22'b1111111111111110001000, 22'b1111111111111000111011, 22'b0000000000000011101110, 22'b1111111111111101011111, 22'b1111111111111011101100, 22'b1111111111111010010011, 22'b1111111111111001010001, 22'b1111111111111111010010, 22'b1111111111110110011110, 22'b0000000000001010010011, 22'b0000000000000011111100, 22'b0000000000001111111001, 22'b0000000000000010110011, 22'b0000000000000001001011, 22'b1111111111110110101100, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b0000000000000110001100, 22'b0000000000000101101011, 22'b0000000000001001011011, 22'b1111111111111111110011, 22'b1111111111110110100111, 22'b0000000000000000010010, 22'b0000000000000000000000, 22'b0000000000001010010100, 22'b1111111111111001100100, 22'b1111111111101110011000, 22'b0000000000010001111101, 22'b1111111111110110100110, 22'b0000000000100101001111, 22'b1111111111111111010111, 22'b1111111111110100101010}, 
{22'b1111111111101101100011, 22'b1111111111111111111100, 22'b1111111111110010111001, 22'b0000000000000111010111, 22'b0000000000001000011011, 22'b1111111111111100101110, 22'b0000000000010000100010, 22'b1111111111111010100011, 22'b1111111111110000101010, 22'b1111111111110100010000, 22'b1111111111110111111101, 22'b1111111111110000110001, 22'b1111111111111000101011, 22'b0000000000000110010011, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b0000000000011010111101, 22'b1111111111111110100111, 22'b1111111111111111111101, 22'b0000000000001101001010, 22'b0000000000001001010111, 22'b1111111111101101011110, 22'b1111111111110011110000, 22'b0000000000000110000011, 22'b1111111111110010001110, 22'b1111111111111111010101, 22'b1111111111110111101100, 22'b1111111111110101010011, 22'b1111111111110010000011, 22'b0000000000001001101010, 22'b0000000000000111010010, 22'b1111111111111011000000, 22'b1111111111111101101011, 22'b1111111111100000110101, 22'b1111111111111010010110, 22'b0000000000000001100101, 22'b1111111111111011110110, 22'b1111111111110110100000, 22'b1111111111111111111000, 22'b0000000000000011110011, 22'b1111111111111100001100, 22'b1111111111111111111010, 22'b1111111111111110111000, 22'b1111111111101010101111, 22'b0000000000000000000001, 22'b0000000000000000000000, 22'b0000000000001010111000, 22'b1111111111111100000001, 22'b0000000000001101100011, 22'b1111111111111001111001, 22'b0000000000001001001101, 22'b1111111111111111111101, 22'b0000000000000111001110, 22'b1111111111110011011110, 22'b1111111111111111111111, 22'b0000000000010000011000, 22'b0000000000001010000000, 22'b0000000000001001010110, 22'b0000000000000000110011, 22'b1111111111110011001101, 22'b1111111111110110011011, 22'b1111111111101010000010, 22'b1111111111111111111100, 22'b0000000000000011011011}, 
{22'b0000000000001001110111, 22'b0000000000000000000101, 22'b0000000000000100001100, 22'b1111111111111111111111, 22'b0000000000000100111010, 22'b1111111111111011101100, 22'b0000000000000111100000, 22'b0000000000000001010110, 22'b0000000000000100010110, 22'b0000000000001010111000, 22'b1111111111110111100100, 22'b1111111111111111010101, 22'b1111111111111111101111, 22'b1111111111111111101110, 22'b1111111111101010111000, 22'b1111111111110110011110, 22'b0000000000010100001011, 22'b1111111111111111000110, 22'b1111111111111110010101, 22'b0000000000000000000000, 22'b1111111111110011110101, 22'b0000000000000000010010, 22'b0000000000001000000001, 22'b0000000000000001001101, 22'b0000000000000001001011, 22'b0000000000001010110101, 22'b0000000000000000000000, 22'b0000000000000001001101, 22'b0000000000000000000000, 22'b1111111111111110011111, 22'b1111111111111001100100, 22'b1111111111101010101100, 22'b0000000000001000011101, 22'b0000000000001010111110, 22'b1111111111111111000100, 22'b1111111111111000011111, 22'b0000000000000000000000, 22'b1111111111101011000011, 22'b1111111111111110100010, 22'b1111111111111111111001, 22'b0000000000000110010001, 22'b1111111111111011110100, 22'b1111111111111111111111, 22'b0000000000011011000111, 22'b0000000000001110010110, 22'b1111111111111111110011, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b1111111111111000010011, 22'b0000000000000100101101, 22'b0000000000000100100111, 22'b0000000000000101100101, 22'b0000000000000101000010, 22'b0000000000001100011011, 22'b0000000000001011001100, 22'b0000000000010101000110, 22'b1111111111111011100001, 22'b0000000000001100100101, 22'b0000000000000100111000, 22'b1111111111110101100100, 22'b0000000000000011100011, 22'b1111111111110011100100, 22'b1111111111110001111011, 22'b1111111111110000000010}, 
{22'b0000000000000000000000, 22'b0000000000000111010011, 22'b1111111111111001110001, 22'b0000000000000000000000, 22'b1111111111111110011011, 22'b1111111111111110111010, 22'b1111111111101010110111, 22'b1111111111111111111111, 22'b0000000000001000000111, 22'b0000000000000111111111, 22'b0000000000000111100110, 22'b1111111111110011010000, 22'b1111111111111101001001, 22'b0000000000001001000101, 22'b1111111111111111111111, 22'b0000000000000000001001, 22'b1111111111100101000100, 22'b1111111111111111111111, 22'b0000000000001011111010, 22'b0000000000000010010000, 22'b0000000000000111100111, 22'b1111111111111100010011, 22'b0000000000000111111111, 22'b0000000000001100111101, 22'b1111111111110100101000, 22'b1111111111110111000011, 22'b1111111111111111110101, 22'b1111111111111101011010, 22'b0000000000000010001001, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b0000000000001010000011, 22'b1111111111101000000000, 22'b0000000000001011100100, 22'b0000000000010000000010, 22'b0000000000000011101110, 22'b0000000000000011100110, 22'b1111111111111100100010, 22'b0000000000000011101011, 22'b1111111111111100100101, 22'b1111111111110111111101, 22'b1111111111111110011000, 22'b0000000000000101010000, 22'b0000000000010110011000, 22'b1111111111100100111000, 22'b1111111111110001101111, 22'b0000000000000110001001, 22'b1111111111111100110111, 22'b0000000000001110011010, 22'b1111111111111000011100, 22'b1111111111110101011010, 22'b1111111111110111000010, 22'b1111111111111111111111, 22'b0000000000000011110110, 22'b1111111111111010111101, 22'b1111111111100101001110, 22'b1111111111111011011011, 22'b1111111111111111101011, 22'b0000000000000001011001, 22'b1111111111101100011110, 22'b0000000000100011110101, 22'b1111111111101110100101, 22'b0000000000010001010101, 22'b0000000000000100111001}, 
{22'b0000000000000010100000, 22'b1111111111111001110111, 22'b0000000000010100000110, 22'b1111111111110110010100, 22'b1111111111110001001011, 22'b0000000000000010111000, 22'b0000000000001001111001, 22'b0000000000001001100111, 22'b1111111111111010010100, 22'b1111111111111010110111, 22'b0000000000000001101011, 22'b0000000000000111010101, 22'b0000000000000111100001, 22'b0000000000000001100110, 22'b1111111111111001011101, 22'b0000000000000100000111, 22'b0000000000001111000100, 22'b1111111111111111101001, 22'b1111111111110111000011, 22'b0000000000000000000000, 22'b0000000000000010011000, 22'b0000000000000000101001, 22'b1111111111110110100111, 22'b0000000000000011100111, 22'b0000000000011001001011, 22'b0000000000000000010100, 22'b0000000000000101110001, 22'b1111111111100110100111, 22'b1111111111111101101011, 22'b0000000000000000010011, 22'b1111111111111001101110, 22'b1111111111110110000001, 22'b0000000000001110101010, 22'b1111111111111111001001, 22'b1111111111111110110010, 22'b1111111111110110001111, 22'b0000000000000100011011, 22'b0000000000001001010110, 22'b1111111111111111101100, 22'b1111111111111110100111, 22'b1111111111111010000001, 22'b0000000000000111010011, 22'b0000000000000000000000, 22'b1111111111101010000010, 22'b0000000000001001111101, 22'b0000000000001100110001, 22'b1111111111111111111111, 22'b0000000000000000110100, 22'b1111111111110010000111, 22'b1111111111111101100110, 22'b1111111111111111111111, 22'b1111111111110101110101, 22'b0000000000000000000000, 22'b1111111111111010011110, 22'b0000000000000001110101, 22'b1111111111100101110110, 22'b1111111111111111111111, 22'b1111111111111111111110, 22'b0000000000001000110011, 22'b0000000000010010000001, 22'b1111111111101001110000, 22'b0000000000010000101001, 22'b0000000000000001001011, 22'b1111111111111101100111}, 
{22'b0000000000001001001101, 22'b0000000000100111101100, 22'b0000000000001111110110, 22'b0000000000001001001000, 22'b1111111111110000101101, 22'b1111111111110101110101, 22'b1111111110101100110100, 22'b1111111111110001011000, 22'b0000000000001100111001, 22'b1111111111111111111111, 22'b0000000000001001011010, 22'b0000000000011011100111, 22'b0000000000000010001110, 22'b0000000000000000001011, 22'b1111111111111111011101, 22'b0000000000000000000000, 22'b1111111111111001111100, 22'b1111111111111001100001, 22'b0000000000000111010111, 22'b1111111111101111111011, 22'b1111111111101010101110, 22'b1111111111111100101101, 22'b1111111111101101010100, 22'b0000000000000000111100, 22'b1111111110110111001001, 22'b0000000000011010000101, 22'b0000000000011111101001, 22'b0000000000010011010100, 22'b1111111111001000001101, 22'b1111111111110101111111, 22'b1111111111101001111111, 22'b1111111111100101000000, 22'b1111111110101111001100, 22'b0000000000010101101001, 22'b1111111111111110100110, 22'b0000000000001010001100, 22'b0000000000000000110000, 22'b1111111111010010001001, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b0000000000000001000001, 22'b0000000000100000100111, 22'b1111111111111001011100, 22'b1111111111101011010111, 22'b0000000000011100101101, 22'b1111111111110001110011, 22'b1111111111110101100111, 22'b1111111111110011011100, 22'b0000000000001111010001, 22'b0000000000010001000000, 22'b1111111111111101110100, 22'b1111111111110100110101, 22'b1111111111111111111011, 22'b1111111111111100011001, 22'b0000000000000000000000, 22'b1111111111110011111011, 22'b0000000000010011011010, 22'b0000000000100010101100, 22'b0000000000010110110001, 22'b1111111111100010111010, 22'b1111111110001001100000, 22'b0000000000011100010101, 22'b0000000000000010111101, 22'b0000000000001010001001}, 
{22'b1111111111111000010001, 22'b0000000000001010110010, 22'b0000000000001010001010, 22'b1111111111111111111100, 22'b1111111111110100000110, 22'b1111111111111101001000, 22'b1111111111110011101110, 22'b1111111111111110001110, 22'b0000000000000100110001, 22'b1111111111111101100110, 22'b1111111111111111000000, 22'b1111111111111110101111, 22'b1111111111111111111110, 22'b1111111111111010001000, 22'b1111111111111111001001, 22'b1111111111111100110010, 22'b0000000000001010000001, 22'b1111111111111111111111, 22'b1111111111101011011111, 22'b0000000000001110111000, 22'b0000000000010011000011, 22'b0000000000001101010001, 22'b1111111111110101110110, 22'b1111111111111011100111, 22'b1111111111110100111011, 22'b1111111111110110101110, 22'b0000000000000111010000, 22'b0000000000000111011111, 22'b0000000000000111001111, 22'b0000000000001011100000, 22'b0000000000000001000110, 22'b0000000000001100010110, 22'b1111111111111110101010, 22'b0000000000000000001001, 22'b0000000000001001101111, 22'b0000000000000100001101, 22'b1111111111111101111000, 22'b1111111111111111101100, 22'b0000000000000000000000, 22'b1111111111110110101000, 22'b1111111111111000110110, 22'b1111111111111100011110, 22'b1111111111110100100000, 22'b0000000000001110011001, 22'b0000000000000000000000, 22'b1111111111111111110100, 22'b1111111111111101010110, 22'b1111111111111011010001, 22'b1111111111100110001110, 22'b1111111111111110110000, 22'b1111111111111000110100, 22'b1111111111111011011101, 22'b1111111111111100110011, 22'b0000000000001000011101, 22'b0000000000010101110100, 22'b0000000000000101111111, 22'b1111111111111111100100, 22'b1111111111110101000001, 22'b1111111111111111000011, 22'b0000000000000000000000, 22'b0000000000001010011010, 22'b1111111111111111010100, 22'b0000000000000001011101, 22'b0000000000000000000000}
};

localparam logic signed [21:0] bias [64] = '{
22'b1111111111111110110011,  // -0.037350185215473175
22'b0000000000001000110000,  // 0.27355897426605225
22'b1111111111111100000010,  // -0.12378914654254913
22'b1111111111111101111011,  // -0.064457006752491
22'b0000000000000001101111,  // 0.05452875792980194
22'b0000000000000011101111,  // 0.11671770364046097
22'b0000000000000100010111,  // 0.13640816509723663
22'b0000000000000010011001,  // 0.07482525706291199
22'b0000000000000001011111,  // 0.04674031585454941
22'b1111111111111001100011,  // -0.20146161317825317
22'b1111111111111100110101,  // -0.09910125285387039
22'b0000000000000100110101,  // 0.15104414522647858
22'b1111111111111100101110,  // -0.10221704095602036
22'b1111111111111011010100,  // -0.1461549550294876
22'b1111111111111101001111,  // -0.08641516417264938
22'b0000000000000101010100,  // 0.16613510251045227
22'b1111111111111101010100,  // -0.0836295336484909
22'b1111111111111110001010,  // -0.05756539851427078
22'b1111111111111110111101,  // -0.03229188174009323
22'b1111111111111111000101,  // -0.028388574719429016
22'b0000000000000100000010,  // 0.1260243058204651
22'b1111111111111110110100,  // -0.037064336240291595
22'b0000000000000110001100,  // 0.19336333870887756
22'b0000000000000000101011,  // 0.02124214917421341
22'b0000000000001111111101,  // 0.4985624849796295
22'b0000000000000000100000,  // 0.0158411655575037
22'b1111111111111101010110,  // -0.08296407759189606
22'b0000000000000011100010,  // 0.11056788265705109
22'b0000000000000000011000,  // 0.01173810102045536
22'b1111111111111100100001,  // -0.10843746364116669
22'b0000000000001000110001,  // 0.27439257502555847
22'b0000000000000010111100,  // 0.09199801832437515
22'b0000000000001000110001,  // 0.27419957518577576
22'b0000000000001000101010,  // 0.27063727378845215
22'b1111111111111000000011,  // -0.24828937649726868
22'b0000000000000010100000,  // 0.07818280160427094
22'b1111111111111111110100,  // -0.005749030504375696
22'b0000000000000011011110,  // 0.10850494354963303
22'b0000000000000100010110,  // 0.13591453433036804
22'b1111111111111100001000,  // -0.12088628858327866
22'b1111111111111110001011,  // -0.05666546896100044
22'b0000000000000010111110,  // 0.09311636537313461
22'b0000000000000001110000,  // 0.05477767437696457
22'b0000000000000000111100,  // 0.029585206881165504
22'b1111111111110110000000,  // -0.31209176778793335
22'b1111111111111101010010,  // -0.08465463668107986
22'b1111111111111010101000,  // -0.16775836050510406
22'b0000000000000100101110,  // 0.14762157201766968
22'b1111111111111000011100,  // -0.23618532717227936
22'b0000000000000010000101,  // 0.06535740196704865
22'b1111111111111011111000,  // -0.12853026390075684
22'b1111111111111011100101,  // -0.13802281022071838
22'b1111111111111011001001,  // -0.15156887471675873
22'b0000000000000010100011,  // 0.07979883998632431
22'b0000000000000101110011,  // 0.18141601979732513
22'b1111111111111110010001,  // -0.054039113223552704
22'b1111111111111111101011,  // -0.010052933357656002
22'b0000000000000010000111,  // 0.06611225008964539
22'b0000000000000001100111,  // 0.05053366720676422
22'b0000000000000000110111,  // 0.026860840618610382
22'b0000000000000001000011,  // 0.03283466026186943
22'b0000000000000100111110,  // 0.15558314323425293
22'b1111111111110110110101,  // -0.2863388657569885
22'b1111111111111101001100   // -0.08769102394580841
};
endpackage