// Width: 26
// NFRAC: 13
package dense_1_26_13;

localparam logic signed [25:0] weights [16][64] = '{ 
{26'b00000000000000100000101001, 26'b11111111111110101100100100, 26'b11111111111111101000110111, 26'b11111111111111100011000000, 26'b11111111111111001100001010, 26'b00000000000000001110001000, 26'b11111111111101111011010000, 26'b00000000000000000000000000, 26'b00000000000000000111011011, 26'b00000000000000100001101110, 26'b00000000000000000000011000, 26'b11111111111111001100001101, 26'b11111111111111111111110111, 26'b00000000000000011010110000, 26'b00000000000000000100010010, 26'b11111111111111011110100000, 26'b00000000000000011101110011, 26'b00000000000000000111100000, 26'b00000000000000000000000000, 26'b11111111111111111111111110, 26'b00000000000000110000001111, 26'b11111111111111010101100100, 26'b11111111111111111101001011, 26'b00000000000000111100100000, 26'b11111111111111010110110110, 26'b11111111111110101000101000, 26'b11111111111111011100101111, 26'b11111111111111100111000000, 26'b11111111111111110010100111, 26'b11111111111111111111110001, 26'b00000000000000000100110101, 26'b00000000000000011111011010, 26'b00000000000000011001000011, 26'b11111111111111111110010100, 26'b00000000000000000000000001, 26'b00000000000000100111110111, 26'b11111111111111111101101100, 26'b11111111111111011111110110, 26'b00000000000000000011011111, 26'b00000000000000011000101001, 26'b11111111111111111110011101, 26'b00000000000000100011001110, 26'b11111111111111011101111001, 26'b00000000000001110110111000, 26'b11111111111111111111110111, 26'b00000000000000111001111011, 26'b00000000000000000000000000, 26'b00000000000000010111100110, 26'b00000000000000011001000110, 26'b11111111111111111100111111, 26'b00000000000000000000000000, 26'b00000000000000010100100010, 26'b00000000000000011011101000, 26'b00000000000000001001111101, 26'b11111111111111110001001111, 26'b11111111111111011000010001, 26'b00000000000001000100101010, 26'b11111111111111000000000011, 26'b00000000000000111011110111, 26'b11111111111111010010101001, 26'b00000000000001100101100001, 26'b11111111111111111111000011, 26'b00000000000000000001011101, 26'b00000000000000001010011000}, 
{26'b00000000000000000000010111, 26'b11111111111111010110111100, 26'b11111111111111101111000011, 26'b11111111111111011100001101, 26'b11111111111111010111010111, 26'b00000000000000001101101001, 26'b11111111111110011111011011, 26'b11111111111111111111101101, 26'b11111111111111100010111010, 26'b00000000000000010110000100, 26'b00000000000000000000110110, 26'b11111111111111110100111110, 26'b00000000000000011001001110, 26'b00000000000000000000000000, 26'b11111111111111111111111110, 26'b00000000000000011010100100, 26'b11111111111111111111001110, 26'b00000000000000000000000010, 26'b11111111111111101000101011, 26'b11111111111111011111111110, 26'b00000000000000111000100111, 26'b11111111111111110101101001, 26'b00000000000000000110001000, 26'b00000000000001011001011101, 26'b00000000000000100000111101, 26'b11111111111111100010100001, 26'b11111111111111100010011100, 26'b11111111111111111111111101, 26'b11111111111111110011000000, 26'b11111111111111001100000111, 26'b11111111111111111000010101, 26'b00000000000000111010001110, 26'b00000000000000100011101010, 26'b00000000000001000110011010, 26'b00000000000001010000100001, 26'b00000000000000000110011101, 26'b11111111111111110000110110, 26'b11111111111111001000011100, 26'b00000000000000000111010000, 26'b00000000000000011000001011, 26'b00000000000000000010111011, 26'b00000000000000011010011011, 26'b11111111111111100100110010, 26'b00000000000000100000010000, 26'b00000000000000010110000011, 26'b00000000000000000110011000, 26'b11111111111111010100011111, 26'b00000000000000001010001011, 26'b00000000000000100001010111, 26'b00000000000000000011110101, 26'b00000000000000000011001011, 26'b00000000000010010100001000, 26'b11111111111111110110011011, 26'b11111111111111110011011101, 26'b11111111111111111001000011, 26'b11111111111111111111000000, 26'b00000000000000100000111000, 26'b11111111111111010000101001, 26'b00000000000001111110000111, 26'b00000000000000000000100111, 26'b00000000000001000010101000, 26'b00000000000000011110101111, 26'b00000000000001101001010011, 26'b00000000000000010010000011}, 
{26'b11111111111111111111000001, 26'b00000000000000000000000000, 26'b11111111111111110101010110, 26'b11111111111111101001011110, 26'b11111111111111101000010111, 26'b00000000000000000101010110, 26'b00000000000010111101100011, 26'b11111111111111111111111111, 26'b11111111111101011101111100, 26'b11111111111111111111111111, 26'b11111111111111111111110001, 26'b11111111111111111101101101, 26'b11111111111111100010111001, 26'b00000000000000000000001010, 26'b11111111111111111110110011, 26'b00000000000000010101100001, 26'b00000000000001110011111001, 26'b11111111111111111111111111, 26'b00000000000000001001001111, 26'b00000000000000000000000010, 26'b00000000000000110100110000, 26'b11111111111110100011101011, 26'b00000000000001001001111010, 26'b11111111111110100100101001, 26'b00000000000001111001011010, 26'b11111111111111010011101010, 26'b11111111111111100000101010, 26'b11111111111110100100001001, 26'b00000000000010100011000000, 26'b00000000000000100011010011, 26'b00000000000000000001011101, 26'b00000000000001000010010001, 26'b00000000000010000010100111, 26'b11111111111101100111000010, 26'b11111111111111110011110001, 26'b00000000000000000100000101, 26'b11111111111111100010011011, 26'b00000000000001110010110100, 26'b11111111111111111010111101, 26'b00000000000000101000000100, 26'b00000000000000101010101000, 26'b00000000000000101111010100, 26'b11111111111111111111111111, 26'b11111111111111111111111110, 26'b11111111111111111101110010, 26'b00000000000000010100000111, 26'b11111111111111011100001100, 26'b11111111111111101010001101, 26'b11111111111111111101110001, 26'b00000000000000110010010110, 26'b11111111111111101001011110, 26'b00000000000000010011001110, 26'b11111111111111111111111100, 26'b00000000000000010001001011, 26'b11111111111111101001100010, 26'b11111111111111111111111111, 26'b11111111111111011000100010, 26'b11111111111110101010010011, 26'b11111111111111111111101111, 26'b00000000000000000000000000, 26'b00000000000011000101011111, 26'b00000000000000000001101010, 26'b11111111111111111111101010, 26'b11111111111111011000011001}, 
{26'b11111111111111000101010110, 26'b11111111111111010000110100, 26'b11111111111110100111010101, 26'b00000000000000100111011101, 26'b11111111111111010111100100, 26'b11111111111101010011101011, 26'b11111111111111110001010100, 26'b11111111111111011000100100, 26'b00000000000000011100101011, 26'b11111111111111111111111111, 26'b00000000000010100001111110, 26'b11111111111111110010011111, 26'b11111111111110011011110110, 26'b00000000000001001010001001, 26'b00000000000000000011001110, 26'b11111111111111111111110011, 26'b11111111111111000111001100, 26'b11111111111111111111111111, 26'b00000000000000000000000000, 26'b11111111111111100011000011, 26'b11111111111101101100101011, 26'b11111111111111110001101101, 26'b11111111111110100110100111, 26'b00000000000000011001011001, 26'b11111111111111001110011111, 26'b11111111111110001010001010, 26'b00000000000000101000000010, 26'b00000000000001011110010010, 26'b00000000000010100101110010, 26'b11111111111111000101001000, 26'b11111111111110110101011011, 26'b00000000000000001001011101, 26'b00000000000001000000000001, 26'b11111111111110010100010100, 26'b11111111111111010111110000, 26'b00000000000000000000000000, 26'b11111111111110100011000100, 26'b00000000000000011111000010, 26'b11111111111111000111100010, 26'b00000000000000001111010001, 26'b00000000000000111010101100, 26'b00000000000000010100000100, 26'b00000000000000000000000000, 26'b00000000000000000010100110, 26'b00000000000001000110101110, 26'b11111111111111100110011010, 26'b11111111111111111111111111, 26'b11111111111111010011111110, 26'b11111111111111111111111111, 26'b11111111111111110011100111, 26'b11111111111110110001001110, 26'b00000000000000001011000111, 26'b11111111111111111111111111, 26'b00000000000000011011111011, 26'b00000000000000101000010111, 26'b00000000000001010010110101, 26'b11111111111110000100001001, 26'b11111111111110001001000111, 26'b11111111111110100101101111, 26'b00000000000001101110111000, 26'b00000000000011011111111000, 26'b11111111111110001100110110, 26'b11111111111111111001000100, 26'b00000000000000110111100101}, 
{26'b00000000000000101011110011, 26'b11111111111110110000110101, 26'b11111111111111011110110011, 26'b11111111111111111111111111, 26'b11111111111111101100010010, 26'b00000000000000101011100011, 26'b00000000000000011000010000, 26'b11111111111111111111111110, 26'b11111111111110110011100010, 26'b11111111111111100001000011, 26'b11111111111111010000110011, 26'b00000000000000000110110001, 26'b00000000000000000000001010, 26'b00000000000000000000000000, 26'b11111111111111111010110100, 26'b00000000000000101101110001, 26'b00000000000000010001000110, 26'b11111111111111001101101101, 26'b00000000000000000011111011, 26'b00000000000000000001101110, 26'b00000000000000011010111001, 26'b11111111111111110000111001, 26'b00000000000000001001100001, 26'b11111111111111111101100011, 26'b00000000000010001000011011, 26'b11111111111111101000001001, 26'b11111111111111011100000000, 26'b11111111111111001100010101, 26'b00000000000000000000000000, 26'b00000000000000010101000101, 26'b00000000000000001110111000, 26'b00000000000000100011000001, 26'b11111111111111111110011010, 26'b00000000000000001001011111, 26'b00000000000000010000101110, 26'b11111111111111111111111111, 26'b00000000000000000000110010, 26'b00000000000001110000110101, 26'b11111111111111011011000001, 26'b11111111111111110110001100, 26'b00000000000000110111011101, 26'b00000000000000011111110110, 26'b11111111111111000001011010, 26'b00000000000000000000110000, 26'b11111111111101110111010000, 26'b11111111111111111111111111, 26'b11111111111111110000010100, 26'b00000000000000000001100001, 26'b11111111111111111111111110, 26'b11111111111111111100111111, 26'b11111111111111111111111111, 26'b00000000000000011000000100, 26'b11111111111111111111010110, 26'b00000000000000101000101011, 26'b11111111111111100111100010, 26'b11111111111110100001111001, 26'b11111111111111000100010011, 26'b11111111111110111110110011, 26'b11111111111110110001011011, 26'b00000000000001011111100110, 26'b00000000000010101111110100, 26'b00000000000001100101011111, 26'b00000000000000001111101100, 26'b11111111111111111111111110}, 
{26'b11111111111111000110111101, 26'b11111111111110101111010010, 26'b00000000000000000000000001, 26'b00000000000000100111010100, 26'b00000000000000100100100001, 26'b11111111111111100100110110, 26'b00000000000001001010100001, 26'b11111111111111111111111111, 26'b00000000000000011111001100, 26'b11111111111111111111111111, 26'b11111111111111111110110011, 26'b11111111111111110110101101, 26'b11111111111111101001011010, 26'b00000000000001001010000000, 26'b11111111111111110100100100, 26'b00000000000000000000000001, 26'b11111111111110110000000001, 26'b11111111111111010010101000, 26'b00000000000000000000000001, 26'b11111111111111111111111111, 26'b11111111111111111001111010, 26'b11111111111111010111110101, 26'b11111111111111010111001100, 26'b00000000000000111011100100, 26'b11111111111111010111010010, 26'b11111111111111111111111000, 26'b00000000000000100000110010, 26'b11111111111111110110101001, 26'b11111111111110001000100110, 26'b11111111111111111111111111, 26'b11111111111111110111011100, 26'b11111111111111111110101011, 26'b11111111111111111110100001, 26'b00000000000000000101001111, 26'b00000000000000010000111000, 26'b00000000000000101100010000, 26'b00000000000000000001101111, 26'b11111111111111110011011100, 26'b11111111111111011110011000, 26'b11111111111111111111110000, 26'b11111111111111101010010111, 26'b11111111111110111100111100, 26'b00000000000000110011001111, 26'b00000000000000000001011000, 26'b00000000000001001101001110, 26'b00000000000000000000000000, 26'b11111111111111111111111110, 26'b00000000000000001100001010, 26'b11111111111111001010010110, 26'b00000000000000011101111101, 26'b00000000000000000000000000, 26'b11111111111111110011000100, 26'b11111111111111010001101111, 26'b00000000000000110001011110, 26'b11111111111111111111111111, 26'b00000000000000101100011011, 26'b00000000000000011011101110, 26'b00000000000000011010000110, 26'b11111111111111111101100111, 26'b11111111111111111110111100, 26'b11111111111110011000100010, 26'b11111111111111101111110110, 26'b11111111111111111000101100, 26'b11111111111111111111111100}, 
{26'b11111111111111011011110011, 26'b11111111111111010101000110, 26'b11111111111111001000110000, 26'b11111111111111110111000110, 26'b11111111111111101110111100, 26'b00000000000000001101010110, 26'b11111111111110100110101000, 26'b11111111111111101100110010, 26'b11111111111111100011010010, 26'b11111111111111111111111110, 26'b11111111111111011011001101, 26'b00000000000000101100100010, 26'b00000000000000000100100011, 26'b00000000000000010001101000, 26'b00000000000000100111111011, 26'b00000000000000000000000010, 26'b00000000000001100110000010, 26'b00000000000000001011011100, 26'b00000000000000011111000101, 26'b00000000000000100010010111, 26'b11111111111111101011111100, 26'b00000000000000101110100000, 26'b11111111111111100000111100, 26'b11111111111110111111110000, 26'b00000000000000010110001100, 26'b00000000000001000010001001, 26'b11111111111111111111011101, 26'b00000000000000000110111001, 26'b11111111111110000110010010, 26'b00000000000000100100101011, 26'b00000000000000100010001100, 26'b11111111111111010000001110, 26'b00000000000000111100010110, 26'b00000000000001010101000101, 26'b00000000000000000000000000, 26'b00000000000000101011110100, 26'b11111111111111111111111111, 26'b00000000000000100100011000, 26'b00000000000000011001011111, 26'b00000000000000000000000000, 26'b11111111111111110000111010, 26'b11111111111111010001011101, 26'b00000000000000010010010111, 26'b00000000000000111101110111, 26'b00000000000001000010011100, 26'b11111111111111101010011110, 26'b11111111111111110101010100, 26'b11111111111111100111101100, 26'b11111111111111101110101100, 26'b00000000000000001111001001, 26'b00000000000000000000011010, 26'b00000000000000000100010111, 26'b00000000000000000000000000, 26'b00000000000000010111001101, 26'b11111111111111101001101010, 26'b00000000000001100010101011, 26'b00000000000000101101100100, 26'b11111111111111111100110101, 26'b00000000000000110001111101, 26'b00000000000000011011110010, 26'b11111111111100101111111111, 26'b11111111111110110110001111, 26'b11111111111111101001111101, 26'b11111111111111111110101110}, 
{26'b00000000000000000000101010, 26'b00000000000000011110100111, 26'b11111111111111111111111101, 26'b11111111111111111111111011, 26'b11111111111111010110110000, 26'b11111111111111111100000000, 26'b11111111111111011111000011, 26'b00000000000000000000000000, 26'b00000000000000000011100001, 26'b00000000000000110001110001, 26'b00000000000000000001110111, 26'b11111111111111001111101000, 26'b11111111111111110111111111, 26'b00000000000000000000000001, 26'b11111111111111111001010000, 26'b11111111111111000110011100, 26'b11111111111110010011011001, 26'b11111111111111111111111101, 26'b11111111111110110010101001, 26'b11111111111111000110111011, 26'b11111111111111001110001001, 26'b00000000000000101100011100, 26'b00000000000000000110000000, 26'b11111111111111101101110001, 26'b11111111111111001000000100, 26'b00000000000000010011111001, 26'b00000000000000000000000000, 26'b00000000000000111111111010, 26'b00000000000001100111001010, 26'b11111111111111111010110110, 26'b00000000000000000000000101, 26'b00000000000000011101100000, 26'b11111111111110101000101011, 26'b11111111111111010000100001, 26'b00000000000000000111000111, 26'b00000000000000001011110110, 26'b11111111111111011100000101, 26'b00000000000000011110101010, 26'b00000000000000010000111001, 26'b11111111111111101100011100, 26'b11111111111111001010010000, 26'b11111111111111111011010000, 26'b00000000000000000100001100, 26'b11111111111111101010101111, 26'b00000000000000000111001001, 26'b00000000000000011101010110, 26'b11111111111111110000101110, 26'b00000000000000000011000011, 26'b00000000000000000000000000, 26'b11111111111111100100000111, 26'b11111111111111001110010011, 26'b00000000000000110101001111, 26'b00000000000000010000001111, 26'b11111111111111101001001100, 26'b00000000000000010000111101, 26'b11111111111111111000000110, 26'b11111111111111000011010001, 26'b11111111111111101110111100, 26'b11111111111111111001010100, 26'b11111111111111110111000001, 26'b00000000000001101010010010, 26'b00000000000000011000011011, 26'b11111111111111111001110011, 26'b11111111111111111111111101}, 
{26'b00000000000000000001111000, 26'b00000000000001001011000111, 26'b11111111111110110101101011, 26'b11111111111111100010011011, 26'b00000000000000101001010011, 26'b11111111111111100101100111, 26'b00000000000010011011000010, 26'b11111111111111011011001011, 26'b11111111111111111111111110, 26'b00000000000000100101100010, 26'b00000000000000100000100010, 26'b11111111111111111111101011, 26'b11111111111111111001110110, 26'b11111111111111000010010010, 26'b00000000000000100100000001, 26'b00000000000000010100011100, 26'b11111111111111100111001100, 26'b11111111111111111111111111, 26'b00000000000000000000000000, 26'b00000000000000000000000010, 26'b00000000000000100001111101, 26'b11111111111111000101001010, 26'b00000000000000110010001100, 26'b00000000000001001110011100, 26'b11111111111111110100110101, 26'b11111111111111111111111101, 26'b11111111111111111101111010, 26'b11111111111111111111111110, 26'b00000000000001011110001110, 26'b00000000000000000000101000, 26'b11111111111111011101000001, 26'b00000000000000000000000000, 26'b00000000000000110001001011, 26'b11111111111110011000001100, 26'b11111111111110111010110010, 26'b00000000000000011001011100, 26'b00000000000000010001101110, 26'b11111111111110110110110110, 26'b11111111111111100111110010, 26'b11111111111111100100100101, 26'b00000000000000110011010101, 26'b00000000000000110010000010, 26'b00000000000000000000000000, 26'b11111111111111011101011100, 26'b00000000000000000000000110, 26'b00000000000000110010100111, 26'b11111111111111111000011101, 26'b11111111111111111111111110, 26'b00000000000000000001011110, 26'b00000000000000011111010111, 26'b11111111111111111000101001, 26'b11111111111111100111001110, 26'b00000000000000101100000011, 26'b11111111111111100100011110, 26'b00000000000000100011110011, 26'b00000000000001001010110101, 26'b00000000000000000101000111, 26'b00000000000000100001101111, 26'b11111111111111001100110001, 26'b11111111111111010001000010, 26'b00000000000001101010011110, 26'b11111111111111101111100001, 26'b00000000000000000101111000, 26'b11111111111111110100000010}, 
{26'b00000000000000000010000100, 26'b11111111111111000110000101, 26'b00000000000000101111001101, 26'b11111111111111011011101010, 26'b11111111111111111111100111, 26'b00000000000000011011000100, 26'b11111111111110110101100000, 26'b00000000000000011000100000, 26'b00000000000000111110110010, 26'b00000000000000010011101111, 26'b00000000000000101110011000, 26'b00000000000000101001010010, 26'b11111111111111011000111111, 26'b11111111111111110110010010, 26'b11111111111111111001011010, 26'b00000000000000000000001001, 26'b11111111111110000101001010, 26'b00000000000000101001010111, 26'b11111111111111111011010111, 26'b00000000000000000011111110, 26'b11111111111111010010111000, 26'b00000000000000001000111100, 26'b00000000000000010011100110, 26'b11111111111111111111111101, 26'b11111111111111000101000101, 26'b11111111111111111001111000, 26'b11111111111111110101100000, 26'b00000000000010011111101110, 26'b11111111111110101011001100, 26'b00000000000000001000100000, 26'b00000000000000001100011010, 26'b11111111111111111000100001, 26'b11111111111111100011101110, 26'b00000000000000001110111010, 26'b11111111111111110101111111, 26'b11111111111111101110110011, 26'b11111111111111101001001101, 26'b11111111111111100101000111, 26'b11111111111111111101001011, 26'b11111111111111011001111011, 26'b00000000000000101001001100, 26'b00000000000000001111110011, 26'b00000000000000111111100101, 26'b00000000000000001011001110, 26'b00000000000000000100101110, 26'b11111111111111011010110001, 26'b00000000000000000000000000, 26'b11111111111111111111111110, 26'b11111111111111111111111100, 26'b00000000000000011000110011, 26'b00000000000000010110101101, 26'b00000000000000100101101111, 26'b11111111111111111111001110, 26'b11111111111111011010011100, 26'b00000000000000000001001001, 26'b00000000000000000000000000, 26'b00000000000000101001010001, 26'b11111111111111100110010010, 26'b11111111111110111001100010, 26'b00000000000001000111110110, 26'b11111111111111011010011000, 26'b00000000000010010100111110, 26'b11111111111111111101011101, 26'b11111111111111010010101000}, 
{26'b11111111111110110110001111, 26'b11111111111111111111110000, 26'b11111111111111001011100100, 26'b00000000000000011101011111, 26'b00000000000000100001101101, 26'b11111111111111110010111001, 26'b00000000000001000010001011, 26'b11111111111111101010001100, 26'b11111111111111000010101001, 26'b11111111111111010001000010, 26'b11111111111111011111110110, 26'b11111111111111000011000101, 26'b11111111111111100010101100, 26'b00000000000000011001001101, 26'b00000000000000000000000000, 26'b00000000000000000000000010, 26'b00000000000001101011110110, 26'b11111111111111111010011110, 26'b11111111111111111111110111, 26'b00000000000000110100101000, 26'b00000000000000100101011110, 26'b11111111111110110101111011, 26'b11111111111111001111000011, 26'b00000000000000011000001100, 26'b11111111111111001000111000, 26'b11111111111111111101010100, 26'b11111111111111011110110001, 26'b11111111111111010101001110, 26'b11111111111111001000001111, 26'b00000000000000100110101011, 26'b00000000000000011101001010, 26'b11111111111111101100000010, 26'b11111111111111110110101100, 26'b11111111111110000011010101, 26'b11111111111111101001011000, 26'b00000000000000000110010101, 26'b11111111111111101111011010, 26'b11111111111111011010000011, 26'b11111111111111111111100010, 26'b00000000000000001111001110, 26'b11111111111111110000110000, 26'b11111111111111111111101010, 26'b11111111111111111011100001, 26'b11111111111110101010111111, 26'b00000000000000000000000110, 26'b00000000000000000000000000, 26'b00000000000000101011100010, 26'b11111111111111110000000101, 26'b00000000000000110110001110, 26'b11111111111111100111100111, 26'b00000000000000100100110111, 26'b11111111111111111111110100, 26'b00000000000000011100111001, 26'b11111111111111001101111010, 26'b11111111111111111111111111, 26'b00000000000001000001100010, 26'b00000000000000101000000001, 26'b00000000000000100101011000, 26'b00000000000000000011001111, 26'b11111111111111001100110100, 26'b11111111111111011001101110, 26'b11111111111110101000001011, 26'b11111111111111111111110000, 26'b00000000000000001101101101}, 
{26'b00000000000000100111011111, 26'b00000000000000000000010101, 26'b00000000000000010000110010, 26'b11111111111111111111111111, 26'b00000000000000010011101001, 26'b11111111111111101110110000, 26'b00000000000000011110000011, 26'b00000000000000000101011011, 26'b00000000000000010001011000, 26'b00000000000000101011100001, 26'b11111111111111011110010001, 26'b11111111111111111101010110, 26'b11111111111111111110111100, 26'b11111111111111111110111000, 26'b11111111111110101011100010, 26'b11111111111111011001111000, 26'b00000000000001010000101101, 26'b11111111111111111100011011, 26'b11111111111111111001010101, 26'b00000000000000000000000010, 26'b11111111111111001111010101, 26'b00000000000000000001001010, 26'b00000000000000100000000111, 26'b00000000000000000100110111, 26'b00000000000000000100101101, 26'b00000000000000101011010100, 26'b00000000000000000000000000, 26'b00000000000000000100110100, 26'b00000000000000000000000000, 26'b11111111111111111001111100, 26'b11111111111111100110010011, 26'b11111111111110101010110001, 26'b00000000000000100001110100, 26'b00000000000000101011111001, 26'b11111111111111111100010000, 26'b11111111111111100001111101, 26'b00000000000000000000000000, 26'b11111111111110101100001101, 26'b11111111111111111010001001, 26'b11111111111111111111100101, 26'b00000000000000011001000101, 26'b11111111111111101111010010, 26'b11111111111111111111111111, 26'b00000000000001101100011101, 26'b00000000000000111001011000, 26'b11111111111111111111001111, 26'b11111111111111111111111101, 26'b11111111111111111111111111, 26'b11111111111111100001001101, 26'b00000000000000010010110100, 26'b00000000000000010010011100, 26'b00000000000000010110010111, 26'b00000000000000010100001001, 26'b00000000000000110001101100, 26'b00000000000000101100110001, 26'b00000000000001010100011010, 26'b11111111111111101110000110, 26'b00000000000000110010010110, 26'b00000000000000010011100011, 26'b11111111111111010110010011, 26'b00000000000000001110001100, 26'b11111111111111001110010010, 26'b11111111111111000111101101, 26'b11111111111111000000001011}, 
{26'b00000000000000000000000010, 26'b00000000000000011101001111, 26'b11111111111111100111000101, 26'b00000000000000000000000000, 26'b11111111111111111001101110, 26'b11111111111111111011101000, 26'b11111111111110101011011101, 26'b11111111111111111111111111, 26'b00000000000000100000011100, 26'b00000000000000011111111110, 26'b00000000000000011110011011, 26'b11111111111111001101000010, 26'b11111111111111110100100101, 26'b00000000000000100100010110, 26'b11111111111111111111111101, 26'b00000000000000000000100111, 26'b11111111111110010100010011, 26'b11111111111111111111111101, 26'b00000000000000101111101011, 26'b00000000000000001001000001, 26'b00000000000000011110011110, 26'b11111111111111110001001111, 26'b00000000000000011111111101, 26'b00000000000000110011110101, 26'b11111111111111010010100001, 26'b11111111111111011100001100, 26'b11111111111111111111010110, 26'b11111111111111110101101010, 26'b00000000000000001000100110, 26'b00000000000000000000000001, 26'b11111111111111111111111111, 26'b00000000000000101000001110, 26'b11111111111110100000000001, 26'b00000000000000101110010000, 26'b00000000000001000000001011, 26'b00000000000000001110111010, 26'b00000000000000001110011001, 26'b11111111111111110010001011, 26'b00000000000000001110101111, 26'b11111111111111110010010101, 26'b11111111111111011111110110, 26'b11111111111111111001100011, 26'b00000000000000010101000011, 26'b00000000000001011001100001, 26'b11111111111110010011100001, 26'b11111111111111000110111100, 26'b00000000000000011000100101, 26'b11111111111111110011011110, 26'b00000000000000111001101011, 26'b11111111111111100001110001, 26'b11111111111111010101101000, 26'b11111111111111011100001000, 26'b11111111111111111111111111, 26'b00000000000000001111011001, 26'b11111111111111101011110111, 26'b11111111111110010100111010, 26'b11111111111111101101101100, 26'b11111111111111111110101100, 26'b00000000000000000101100100, 26'b11111111111110110001111000, 26'b00000000000010001111010111, 26'b11111111111110111010010101, 26'b00000000000001000101010101, 26'b00000000000000010011100111}, 
{26'b00000000000000001010000001, 26'b11111111111111100111011101, 26'b00000000000001010000011010, 26'b11111111111111011001010011, 26'b11111111111111000100101100, 26'b00000000000000001011100000, 26'b00000000000000100111100110, 26'b00000000000000100110011111, 26'b11111111111111101001010010, 26'b11111111111111101011011100, 26'b00000000000000000110101110, 26'b00000000000000011101010100, 26'b00000000000000011110000100, 26'b00000000000000000110011011, 26'b11111111111111100101110111, 26'b00000000000000010000011100, 26'b00000000000000111100010000, 26'b11111111111111111110100100, 26'b11111111111111011100001100, 26'b00000000000000000000000001, 26'b00000000000000001001100001, 26'b00000000000000000010100110, 26'b11111111111111011010011110, 26'b00000000000000001110011101, 26'b00000000000001100100101111, 26'b00000000000000000001010010, 26'b00000000000000010111000111, 26'b11111111111110011010011110, 26'b11111111111111110110101100, 26'b00000000000000000001001100, 26'b11111111111111100110111000, 26'b11111111111111011000000111, 26'b00000000000000111010101010, 26'b11111111111111111100100110, 26'b11111111111111111011001011, 26'b11111111111111011000111100, 26'b00000000000000010001101110, 26'b00000000000000100101011001, 26'b11111111111111111110110001, 26'b11111111111111111010011100, 26'b11111111111111101000000111, 26'b00000000000000011101001110, 26'b00000000000000000000000000, 26'b11111111111110101000001001, 26'b00000000000000100111110101, 26'b00000000000000110011000100, 26'b11111111111111111111111110, 26'b00000000000000000011010000, 26'b11111111111111001000011101, 26'b11111111111111110110011010, 26'b11111111111111111111111111, 26'b11111111111111010111010110, 26'b00000000000000000000000000, 26'b11111111111111101001111001, 26'b00000000000000000111010101, 26'b11111111111110010111011001, 26'b11111111111111111111111111, 26'b11111111111111111111111000, 26'b00000000000000100011001110, 26'b00000000000001001000000100, 26'b11111111111110100111000011, 26'b00000000000001000010100101, 26'b00000000000000000100101111, 26'b11111111111111110110011101}, 
{26'b00000000000000100100110101, 26'b00000000000010011110110000, 26'b00000000000000111111011011, 26'b00000000000000100100100000, 26'b11111111111111000010110111, 26'b11111111111111010111010111, 26'b11111111111010110011010001, 26'b11111111111111000101100000, 26'b00000000000000110011100101, 26'b11111111111111111111111111, 26'b00000000000000100101101001, 26'b00000000000001101110011111, 26'b00000000000000001000111001, 26'b00000000000000000000101101, 26'b11111111111111111101110101, 26'b00000000000000000000000001, 26'b11111111111111100111110000, 26'b11111111111111100110000100, 26'b00000000000000011101011101, 26'b11111111111110111111101111, 26'b11111111111110101010111000, 26'b11111111111111110010110111, 26'b11111111111110110101010000, 26'b00000000000000000011110001, 26'b11111111111011011100100110, 26'b00000000000001101000010111, 26'b00000000000001111110100111, 26'b00000000000001001101010000, 26'b11111111111100100000110110, 26'b11111111111111010111111101, 26'b11111111111110100111111100, 26'b11111111111110010100000001, 26'b11111111111010111100110010, 26'b00000000000001010110100101, 26'b11111111111111111010011001, 26'b00000000000000101000110011, 26'b00000000000000000011000010, 26'b11111111111101001000100101, 26'b00000000000000000000000010, 26'b00000000000000000000000000, 26'b00000000000000000100000101, 26'b00000000000010000010011110, 26'b11111111111111100101110000, 26'b11111111111110101101011101, 26'b00000000000001110010110111, 26'b11111111111111000111001100, 26'b11111111111111010110011110, 26'b11111111111111001101110000, 26'b00000000000000111101000111, 26'b00000000000001000100000000, 26'b11111111111111110111010011, 26'b11111111111111010011010100, 26'b11111111111111111111101110, 26'b11111111111111110001100111, 26'b00000000000000000000000000, 26'b11111111111111001111101110, 26'b00000000000001001101101000, 26'b00000000000010001010110010, 26'b00000000000001011011000101, 26'b11111111111110001011101010, 26'b11111111111000100110000000, 26'b00000000000001110001010101, 26'b00000000000000001011110101, 26'b00000000000000101000100100}, 
{26'b11111111111111100001000101, 26'b00000000000000101011001011, 26'b00000000000000101000101001, 26'b11111111111111111111110011, 26'b11111111111111010000011001, 26'b11111111111111110100100001, 26'b11111111111111001110111001, 26'b11111111111111111000111000, 26'b00000000000000010011000101, 26'b11111111111111110110011001, 26'b11111111111111111100000010, 26'b11111111111111111010111111, 26'b11111111111111111111111010, 26'b11111111111111101000100010, 26'b11111111111111111100100101, 26'b11111111111111110011001010, 26'b00000000000000101000000111, 26'b11111111111111111111111111, 26'b11111111111110101101111100, 26'b00000000000000111011100001, 26'b00000000000001001100001101, 26'b00000000000000110101000100, 26'b11111111111111010111011010, 26'b11111111111111101110011101, 26'b11111111111111010011101110, 26'b11111111111111011010111001, 26'b00000000000000011101000011, 26'b00000000000000011101111100, 26'b00000000000000011100111100, 26'b00000000000000101110000011, 26'b00000000000000000100011000, 26'b00000000000000110001011010, 26'b11111111111111111010101001, 26'b00000000000000000000100111, 26'b00000000000000100110111111, 26'b00000000000000010000110101, 26'b11111111111111110111100011, 26'b11111111111111111110110010, 26'b00000000000000000000000000, 26'b11111111111111011010100011, 26'b11111111111111100011011010, 26'b11111111111111110001111000, 26'b11111111111111010010000010, 26'b00000000000000111001100100, 26'b00000000000000000000000010, 26'b11111111111111111111010010, 26'b11111111111111110101011011, 26'b11111111111111101101000110, 26'b11111111111110011000111000, 26'b11111111111111111011000010, 26'b11111111111111100011010001, 26'b11111111111111101101110111, 26'b11111111111111110011001101, 26'b00000000000000100001110110, 26'b00000000000001010111010011, 26'b00000000000000010111111111, 26'b11111111111111111110010011, 26'b11111111111111010100000110, 26'b11111111111111111100001111, 26'b00000000000000000000000010, 26'b00000000000000101001101011, 26'b11111111111111111101010010, 26'b00000000000000000101110111, 26'b00000000000000000000000000}
};

localparam logic signed [25:0] bias [64] = '{
26'b11111111111111111011001110,  // -0.037350185215473175
26'b00000000000000100011000000,  // 0.27355897426605225
26'b11111111111111110000001001,  // -0.12378914654254913
26'b11111111111111110111101111,  // -0.064457006752491
26'b00000000000000000110111110,  // 0.05452875792980194
26'b00000000000000001110111100,  // 0.11671770364046097
26'b00000000000000010001011101,  // 0.13640816509723663
26'b00000000000000001001100100,  // 0.07482525706291199
26'b00000000000000000101111110,  // 0.04674031585454941
26'b11111111111111100110001101,  // -0.20146161317825317
26'b11111111111111110011010100,  // -0.09910125285387039
26'b00000000000000010011010101,  // 0.15104414522647858
26'b11111111111111110010111010,  // -0.10221704095602036
26'b11111111111111101101010010,  // -0.1461549550294876
26'b11111111111111110100111100,  // -0.08641516417264938
26'b00000000000000010101010000,  // 0.16613510251045227
26'b11111111111111110101010010,  // -0.0836295336484909
26'b11111111111111111000101000,  // -0.05756539851427078
26'b11111111111111111011110111,  // -0.03229188174009323
26'b11111111111111111100010111,  // -0.028388574719429016
26'b00000000000000010000001000,  // 0.1260243058204651
26'b11111111111111111011010000,  // -0.037064336240291595
26'b00000000000000011000110000,  // 0.19336333870887756
26'b00000000000000000010101110,  // 0.02124214917421341
26'b00000000000000111111110100,  // 0.4985624849796295
26'b00000000000000000010000001,  // 0.0158411655575037
26'b11111111111111110101011000,  // -0.08296407759189606
26'b00000000000000001110001001,  // 0.11056788265705109
26'b00000000000000000001100000,  // 0.01173810102045536
26'b11111111111111110010000111,  // -0.10843746364116669
26'b00000000000000100011000111,  // 0.27439257502555847
26'b00000000000000001011110001,  // 0.09199801832437515
26'b00000000000000100011000110,  // 0.27419957518577576
26'b00000000000000100010101001,  // 0.27063727378845215
26'b11111111111111100000001110,  // -0.24828937649726868
26'b00000000000000001010000000,  // 0.07818280160427094
26'b11111111111111111111010000,  // -0.005749030504375696
26'b00000000000000001101111000,  // 0.10850494354963303
26'b00000000000000010001011001,  // 0.13591453433036804
26'b11111111111111110000100001,  // -0.12088628858327866
26'b11111111111111111000101111,  // -0.05666546896100044
26'b00000000000000001011111010,  // 0.09311636537313461
26'b00000000000000000111000000,  // 0.05477767437696457
26'b00000000000000000011110010,  // 0.029585206881165504
26'b11111111111111011000000011,  // -0.31209176778793335
26'b11111111111111110101001010,  // -0.08465463668107986
26'b11111111111111101010100001,  // -0.16775836050510406
26'b00000000000000010010111001,  // 0.14762157201766968
26'b11111111111111100001110001,  // -0.23618532717227936
26'b00000000000000001000010111,  // 0.06535740196704865
26'b11111111111111101111100011,  // -0.12853026390075684
26'b11111111111111101110010101,  // -0.13802281022071838
26'b11111111111111101100100110,  // -0.15156887471675873
26'b00000000000000001010001101,  // 0.07979883998632431
26'b00000000000000010111001110,  // 0.18141601979732513
26'b11111111111111111001000101,  // -0.054039113223552704
26'b11111111111111111110101101,  // -0.010052933357656002
26'b00000000000000001000011101,  // 0.06611225008964539
26'b00000000000000000110011101,  // 0.05053366720676422
26'b00000000000000000011011100,  // 0.026860840618610382
26'b00000000000000000100001100,  // 0.03283466026186943
26'b00000000000000010011111010,  // 0.15558314323425293
26'b11111111111111011011010110,  // -0.2863388657569885
26'b11111111111111110100110001   // -0.08769102394580841
};
endpackage