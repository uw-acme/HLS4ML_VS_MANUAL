// Width: 13
// NFRAC: 6
package dense_2_13_6;

localparam logic signed [12:0] weights [64][32] = '{ 
{13'b0000000010001, 13'b0000000000000, 13'b1111111110011, 13'b1111111111110, 13'b0000000010000, 13'b0000000000000, 13'b1111111110110, 13'b1111111111111, 13'b1111111101110, 13'b0000000000101, 13'b0000000000000, 13'b1111111111111, 13'b1111111111111, 13'b1111111110011, 13'b1111111111100, 13'b1111111101111, 13'b0000000000000, 13'b1111111111111, 13'b1111111110011, 13'b1111111110101, 13'b0000000000000, 13'b0000000000000, 13'b1111111111111, 13'b1111111111111, 13'b0000000000000, 13'b0000000000110, 13'b0000000011000, 13'b0000000001011, 13'b1111111111111, 13'b0000000000011, 13'b1111111100101, 13'b0000000000000}, 
{13'b1111111111001, 13'b1111111110110, 13'b1111111110111, 13'b1111111111100, 13'b1111111111111, 13'b0000000000010, 13'b1111111110001, 13'b0000000000000, 13'b0000000000000, 13'b1111111111011, 13'b0000000001001, 13'b1111111111101, 13'b1111111111100, 13'b1111111110010, 13'b0000000000000, 13'b1111111111100, 13'b0000000000000, 13'b1111111110011, 13'b0000000001010, 13'b0000000001110, 13'b1111111111101, 13'b1111111111111, 13'b1111111111111, 13'b0000000000001, 13'b1111111111011, 13'b0000000010001, 13'b0000000001111, 13'b0000000000000, 13'b0000000000001, 13'b1111111100000, 13'b0000000000000, 13'b0000000000000}, 
{13'b0000000000100, 13'b1111111111000, 13'b1111111110111, 13'b1111111111101, 13'b1111111111011, 13'b1111111111010, 13'b1111111110100, 13'b0000000000000, 13'b1111111110111, 13'b0000000000000, 13'b0000000000000, 13'b1111111111010, 13'b0000000000101, 13'b1111111111011, 13'b1111111111111, 13'b1111111111101, 13'b0000000000000, 13'b0000000000110, 13'b0000000000011, 13'b0000000001110, 13'b0000000000010, 13'b1111111111010, 13'b0000000000000, 13'b0000000000010, 13'b1111111111110, 13'b0000000001101, 13'b0000000001001, 13'b0000000000110, 13'b1111111111111, 13'b1111111110110, 13'b1111111111111, 13'b0000000000110}, 
{13'b0000000001000, 13'b0000000000001, 13'b0000000000011, 13'b1111111111111, 13'b1111111011111, 13'b0000000000000, 13'b0000000000000, 13'b0000000001110, 13'b0000000001111, 13'b1111111111111, 13'b1111111111111, 13'b0000000000000, 13'b0000000000000, 13'b0000000000000, 13'b1111111111110, 13'b0000000001101, 13'b0000000000000, 13'b1111111111110, 13'b1111111111111, 13'b1111111110100, 13'b1111111111100, 13'b0000000000011, 13'b1111111111011, 13'b1111111111111, 13'b0000000000000, 13'b1111111111100, 13'b0000000000100, 13'b1111111111111, 13'b1111111111111, 13'b1111111111111, 13'b1111111110010, 13'b0000000010011}, 
{13'b1111111010100, 13'b1111111111110, 13'b1111111111111, 13'b0000000000000, 13'b1111111111110, 13'b0000000000000, 13'b1111111111100, 13'b1111111110110, 13'b0000000000011, 13'b1111111111110, 13'b1111111111111, 13'b1111111111111, 13'b1111111111111, 13'b0000000001101, 13'b0000000000000, 13'b0000000010101, 13'b1111111111111, 13'b0000000001101, 13'b1111111100110, 13'b0000000000000, 13'b1111111111000, 13'b0000000001010, 13'b0000000010000, 13'b0000000000000, 13'b0000000000010, 13'b0000000001010, 13'b0000000001111, 13'b0000000000001, 13'b1111111111111, 13'b1111111111111, 13'b1111111111111, 13'b0000000001110}, 
{13'b0000000000011, 13'b1111111111111, 13'b0000000001001, 13'b1111111010110, 13'b1111110100111, 13'b1111111101001, 13'b0000000010110, 13'b1111111011000, 13'b1111111111111, 13'b1111111010100, 13'b1111111011111, 13'b1111111101010, 13'b0000000010110, 13'b1111111111111, 13'b1111111111111, 13'b0000000000000, 13'b1111111111111, 13'b1111111111111, 13'b1111111110111, 13'b1111111111111, 13'b1111111100000, 13'b0000000000000, 13'b0000000001011, 13'b1111111111111, 13'b0000000000001, 13'b0000000010001, 13'b0000000000011, 13'b1111111111111, 13'b1111111111111, 13'b0000000001101, 13'b1111111111101, 13'b0000000001100}, 
{13'b1111111111101, 13'b1111111110101, 13'b1111111110000, 13'b1111111111100, 13'b1111111101101, 13'b0000000000100, 13'b1111111110100, 13'b1111111110110, 13'b1111111100101, 13'b0000000000011, 13'b1111111111111, 13'b1111111110101, 13'b0000000000111, 13'b1111111111111, 13'b1111111111101, 13'b1111111011100, 13'b1111111111111, 13'b0000000000101, 13'b0000000001100, 13'b1111111110101, 13'b1111111110110, 13'b1111111111011, 13'b1111111111111, 13'b0000000000001, 13'b1111111111101, 13'b1111111010110, 13'b1111111101111, 13'b1111111111101, 13'b0000000000000, 13'b1111111111110, 13'b0000000000001, 13'b1111111111111}, 
{13'b1111111110110, 13'b1111111111010, 13'b1111111111010, 13'b1111111110000, 13'b1111111111000, 13'b1111111111111, 13'b0000000000110, 13'b1111111111010, 13'b0000000001100, 13'b0000000000000, 13'b0000000000000, 13'b1111111111111, 13'b0000000001110, 13'b0000000000000, 13'b1111111111111, 13'b1111111111011, 13'b1111111111111, 13'b0000000000000, 13'b1111111111111, 13'b0000000000000, 13'b1111111111111, 13'b1111111111111, 13'b0000000000000, 13'b1111111111111, 13'b0000000000010, 13'b1111111110100, 13'b0000000000000, 13'b1111111111111, 13'b1111111111011, 13'b1111111111111, 13'b0000000000000, 13'b1111111111111}, 
{13'b1111111100001, 13'b1111111111100, 13'b1111111100111, 13'b0000000000111, 13'b0000000011111, 13'b1111111111111, 13'b1111111111110, 13'b0000000001111, 13'b1111111100011, 13'b1111111111101, 13'b0000000000000, 13'b1111111110011, 13'b1111111111111, 13'b0000000000100, 13'b1111111110011, 13'b0000000110000, 13'b1111111111111, 13'b0000000000010, 13'b0000000001101, 13'b0000000001111, 13'b0000000000000, 13'b1111111101010, 13'b0000000000000, 13'b0000000011010, 13'b1111111110100, 13'b0000000101100, 13'b1111111110110, 13'b1111111110010, 13'b1111111100001, 13'b1111111100010, 13'b0000000000000, 13'b0000000000011}, 
{13'b0000000000000, 13'b1111111111111, 13'b1111111111011, 13'b0000000000000, 13'b0000000010011, 13'b1111111111110, 13'b1111111111011, 13'b0000000000101, 13'b0000000000110, 13'b0000000000000, 13'b1111111111111, 13'b1111111111111, 13'b1111111111111, 13'b1111111111000, 13'b1111111111111, 13'b0000000000000, 13'b0000000000000, 13'b1111111111111, 13'b0000000000000, 13'b0000000000101, 13'b0000000000001, 13'b1111111111111, 13'b0000000000000, 13'b0000000000000, 13'b0000000000010, 13'b1111111110111, 13'b0000000000100, 13'b0000000001111, 13'b1111111111111, 13'b0000000000000, 13'b0000000000011, 13'b0000000000100}, 
{13'b0000000000110, 13'b0000000000000, 13'b1111111111001, 13'b1111111101111, 13'b1111111001101, 13'b0000000001000, 13'b0000000000000, 13'b1111111001011, 13'b0000000000010, 13'b1111111111111, 13'b0000000000000, 13'b1111111111111, 13'b0000000000000, 13'b0000000000000, 13'b1111111111110, 13'b1111111100111, 13'b1111111111111, 13'b0000000001110, 13'b0000000001000, 13'b0000000001100, 13'b1111111100011, 13'b1111111101001, 13'b0000000000111, 13'b1111111111101, 13'b1111111111101, 13'b0000000010110, 13'b1111111111001, 13'b1111111111111, 13'b1111111111111, 13'b0000000001101, 13'b1111111111111, 13'b0000000000000}, 
{13'b1111111110011, 13'b1111111100000, 13'b0000000000000, 13'b1111111111111, 13'b0000000010101, 13'b1111111101110, 13'b1111111110001, 13'b0000000000111, 13'b1111111111111, 13'b0000000001001, 13'b0000000000100, 13'b1111111111011, 13'b0000000000000, 13'b0000000000000, 13'b1111111111110, 13'b1111111101111, 13'b0000000001011, 13'b0000000000001, 13'b0000000010011, 13'b0000000000101, 13'b0000000000000, 13'b1111111111101, 13'b0000000001000, 13'b1111111111010, 13'b1111111101100, 13'b1111111111111, 13'b0000000001011, 13'b1111111111111, 13'b0000000000000, 13'b1111111111001, 13'b0000000001000, 13'b0000000010001}, 
{13'b0000000000000, 13'b0000000000000, 13'b0000000001110, 13'b0000000000000, 13'b1111111111101, 13'b0000000001011, 13'b0000000000101, 13'b1111111111111, 13'b0000000000000, 13'b1111111110111, 13'b1111111111100, 13'b1111111110101, 13'b1111111111111, 13'b0000000000011, 13'b1111111111011, 13'b0000000110101, 13'b0000000000000, 13'b1111111111001, 13'b1111111110011, 13'b1111111111111, 13'b0000000001100, 13'b0000000001000, 13'b0000000000000, 13'b1111111111111, 13'b0000000001110, 13'b0000000010001, 13'b0000000011111, 13'b0000000000000, 13'b0000000000000, 13'b0000000000000, 13'b1111111111111, 13'b1111111111011}, 
{13'b1111111110110, 13'b0000000000011, 13'b0000000000010, 13'b1111111110000, 13'b1111111101110, 13'b0000000011110, 13'b0000000000011, 13'b0000000000000, 13'b1111111110101, 13'b1111111111010, 13'b0000000001000, 13'b0000000000100, 13'b0000000000000, 13'b1111111111010, 13'b0000000010010, 13'b1111111111111, 13'b1111111111111, 13'b0000000000000, 13'b0000000000000, 13'b1111111111101, 13'b0000000000101, 13'b0000000000001, 13'b0000000000111, 13'b1111111111111, 13'b0000000000000, 13'b0000000101010, 13'b1111111111100, 13'b1111111111110, 13'b1111111111111, 13'b1111111111001, 13'b1111111111101, 13'b0000000001011}, 
{13'b0000000000011, 13'b0000000000100, 13'b0000000010100, 13'b1111111111101, 13'b0000000000110, 13'b0000000010110, 13'b0000000000000, 13'b1111111111110, 13'b0000000000111, 13'b1111111111000, 13'b1111111111111, 13'b1111111111000, 13'b0000000000000, 13'b0000000011001, 13'b1111111111110, 13'b0000000000000, 13'b0000000001111, 13'b0000000000000, 13'b0000000000000, 13'b1111111101011, 13'b1111111110000, 13'b1111111111101, 13'b1111111111111, 13'b1111111110110, 13'b1111111111101, 13'b1111111111010, 13'b1111111110011, 13'b1111111110010, 13'b0000000000001, 13'b0000000000111, 13'b1111111100110, 13'b0000000000000}, 
{13'b1111111101100, 13'b0000000000000, 13'b1111111111111, 13'b1111111111100, 13'b1111111111111, 13'b0000000001000, 13'b1111111111011, 13'b0000000010001, 13'b1111111101000, 13'b1111111111111, 13'b0000000000000, 13'b1111111111111, 13'b0000000000000, 13'b0000000000000, 13'b1111111111111, 13'b1111111111010, 13'b0000000000101, 13'b0000000001011, 13'b1111111111111, 13'b1111111101111, 13'b1111111111100, 13'b0000000000111, 13'b0000000000100, 13'b0000000000000, 13'b0000000000000, 13'b0000000000101, 13'b1111111110000, 13'b0000000000000, 13'b1111111111111, 13'b0000000000000, 13'b0000000000000, 13'b1111111110111}, 
{13'b1111111101010, 13'b1111111111111, 13'b1111111111111, 13'b1111111111110, 13'b1111111111111, 13'b0000000000110, 13'b0000000000000, 13'b0000000000010, 13'b0000000000010, 13'b0000000000100, 13'b0000000000101, 13'b0000000001010, 13'b0000000000001, 13'b1111111111001, 13'b0000000000000, 13'b0000000011000, 13'b0000000000000, 13'b0000000000000, 13'b1111111111111, 13'b0000000000111, 13'b0000000001001, 13'b0000000000001, 13'b0000000000010, 13'b1111111111110, 13'b1111111111101, 13'b0000000000001, 13'b1111111111011, 13'b1111111110111, 13'b0000000001101, 13'b1111111111110, 13'b0000000000010, 13'b1111111110011}, 
{13'b0000000000000, 13'b1111111111111, 13'b0000000000010, 13'b0000000000000, 13'b0000000111010, 13'b1111111111111, 13'b0000000000000, 13'b1111111111111, 13'b0000000000111, 13'b1111111111011, 13'b0000000000000, 13'b0000000000000, 13'b0000000000000, 13'b0000000001000, 13'b0000000000000, 13'b1111111110110, 13'b1111111111111, 13'b1111111111011, 13'b0000000010100, 13'b0000000000000, 13'b1111111111111, 13'b1111111111111, 13'b0000000000000, 13'b1111111111111, 13'b0000000000000, 13'b0000000000100, 13'b0000000000000, 13'b0000000000000, 13'b1111111111111, 13'b1111111111111, 13'b0000000000000, 13'b0000000000010}, 
{13'b1111111111111, 13'b0000000000001, 13'b1111111111111, 13'b0000000000011, 13'b1111111111101, 13'b1111111111000, 13'b1111111111100, 13'b0000000010001, 13'b0000000000000, 13'b0000000000110, 13'b1111111111111, 13'b0000000000100, 13'b1111111111101, 13'b1111111110101, 13'b1111111110011, 13'b0000000000000, 13'b1111111111111, 13'b1111111111101, 13'b0000000000000, 13'b0000000000000, 13'b1111111111111, 13'b0000000000100, 13'b0000000000010, 13'b1111111110111, 13'b0000000000111, 13'b1111111110101, 13'b0000000000000, 13'b0000000000000, 13'b1111111110101, 13'b0000000000000, 13'b0000000000010, 13'b1111111111110}, 
{13'b1111111111111, 13'b1111111111001, 13'b0000000000000, 13'b1111111111100, 13'b0000000001101, 13'b1111111111111, 13'b1111111111110, 13'b0000000000110, 13'b1111111100110, 13'b0000000000000, 13'b1111111111101, 13'b1111111111111, 13'b0000000010110, 13'b0000000001110, 13'b1111111111001, 13'b1111111111110, 13'b1111111111111, 13'b0000000000000, 13'b1111111111111, 13'b0000000000000, 13'b0000000000000, 13'b1111111110111, 13'b1111111111000, 13'b0000000001000, 13'b0000000000000, 13'b1111111110111, 13'b0000000000001, 13'b1111111111010, 13'b1111111111101, 13'b0000000001000, 13'b0000000000000, 13'b1111111110000}, 
{13'b0000000101000, 13'b0000000010101, 13'b1111111110000, 13'b0000000000000, 13'b1111111101001, 13'b0000000000000, 13'b0000000001110, 13'b0000000000001, 13'b0000000001110, 13'b1111111111111, 13'b1111111110110, 13'b1111111111010, 13'b0000000001001, 13'b0000000000001, 13'b1111111111001, 13'b0000000001000, 13'b0000000100010, 13'b1111111110111, 13'b1111111101101, 13'b0000000000000, 13'b1111111111110, 13'b1111111110100, 13'b1111111111111, 13'b1111111111111, 13'b0000000000101, 13'b1111111101000, 13'b0000000000101, 13'b1111111111111, 13'b0000000000000, 13'b0000000000110, 13'b1111111111110, 13'b0000000000011}, 
{13'b1111111111010, 13'b1111111110011, 13'b1111111111101, 13'b1111111110101, 13'b1111111111110, 13'b0000000000011, 13'b0000000000000, 13'b1111111111111, 13'b0000000000010, 13'b1111111111111, 13'b0000000000000, 13'b1111111110010, 13'b0000000000110, 13'b0000000000101, 13'b1111111111001, 13'b0000000011100, 13'b1111111111111, 13'b0000000000000, 13'b1111111111111, 13'b0000000000000, 13'b0000000010100, 13'b1111111100001, 13'b1111111111001, 13'b1111111111100, 13'b1111111111110, 13'b0000000001100, 13'b1111111111100, 13'b0000000000001, 13'b0000000011110, 13'b1111111011111, 13'b1111111101000, 13'b0000000000001}, 
{13'b0000000000001, 13'b1111111111100, 13'b1111111111111, 13'b0000000000000, 13'b1111111010001, 13'b1111111011001, 13'b0000000000000, 13'b1111111111111, 13'b1111111101111, 13'b0000000000001, 13'b0000000000000, 13'b1111111111110, 13'b0000000000000, 13'b1111111111100, 13'b1111111111100, 13'b1111111111011, 13'b1111111110110, 13'b0000000010010, 13'b0000000000000, 13'b0000000000010, 13'b1111111111111, 13'b1111111111011, 13'b0000000000000, 13'b1111111111010, 13'b0000000001110, 13'b1111111011000, 13'b0000000001110, 13'b1111111111111, 13'b1111111111111, 13'b0000000001100, 13'b1111111111111, 13'b0000000001111}, 
{13'b1111111111111, 13'b0000000000000, 13'b1111111111101, 13'b0000000000100, 13'b0000000000011, 13'b1111111101010, 13'b0000000000000, 13'b0000000000100, 13'b0000000100101, 13'b1111111111111, 13'b0000000000000, 13'b0000000000011, 13'b0000000010110, 13'b1111111111101, 13'b0000000000000, 13'b0000000000110, 13'b1111111111111, 13'b0000000000001, 13'b1111111111111, 13'b0000000000000, 13'b1111111101110, 13'b0000000000010, 13'b0000000000100, 13'b0000000000001, 13'b1111111111111, 13'b0000000001101, 13'b0000000000000, 13'b0000000001000, 13'b1111111100101, 13'b0000000000110, 13'b0000000011001, 13'b0000000000000}, 
{13'b1111111101001, 13'b0000000001101, 13'b1111111101111, 13'b0000000000111, 13'b1111111111001, 13'b0000000000000, 13'b0000000011111, 13'b1111111110001, 13'b1111111101101, 13'b0000000001010, 13'b1111111110001, 13'b1111111111110, 13'b1111111111111, 13'b0000000010110, 13'b1111111111111, 13'b1111111101100, 13'b1111111111111, 13'b0000000011100, 13'b1111111100001, 13'b1111111111110, 13'b0000000010100, 13'b1111111101000, 13'b0000000000011, 13'b1111111111111, 13'b0000000010001, 13'b1111111011111, 13'b1111111101000, 13'b1111111110011, 13'b1111111111111, 13'b0000000000110, 13'b0000000000001, 13'b0000000001011}, 
{13'b1111111111010, 13'b0000000000011, 13'b1111111111111, 13'b0000000001001, 13'b1111111111101, 13'b0000000001110, 13'b0000000000000, 13'b1111111111111, 13'b1111111111111, 13'b0000000000000, 13'b0000000000000, 13'b1111111111111, 13'b1111111111111, 13'b0000000100001, 13'b0000000000000, 13'b0000000001100, 13'b0000000000000, 13'b1111111110010, 13'b1111111111011, 13'b1111111111111, 13'b1111111111110, 13'b0000000000010, 13'b1111111111111, 13'b1111111110100, 13'b1111111111111, 13'b0000000010010, 13'b0000000010011, 13'b1111111111111, 13'b1111111111110, 13'b0000000000000, 13'b1111111111111, 13'b1111111111001}, 
{13'b1111111111010, 13'b0000000000000, 13'b0000000010001, 13'b0000000000000, 13'b0000000000000, 13'b1111111111000, 13'b0000000000000, 13'b1111111001000, 13'b0000000001101, 13'b0000000000000, 13'b0000000000001, 13'b1111111101000, 13'b0000000000000, 13'b1111111110111, 13'b1111111111101, 13'b0000000000000, 13'b0000000000001, 13'b0000000000000, 13'b0000000000111, 13'b0000000000000, 13'b1111111111111, 13'b0000000010101, 13'b0000000011000, 13'b1111111110001, 13'b1111111110110, 13'b0000000001111, 13'b1111111101100, 13'b0000000000001, 13'b1111111111111, 13'b1111111111111, 13'b1111111111111, 13'b0000000001011}, 
{13'b1111111111000, 13'b1111111111111, 13'b1111111110000, 13'b1111111110011, 13'b1111111111111, 13'b1111111110111, 13'b0000000000000, 13'b0000000000101, 13'b1111111110000, 13'b1111111111010, 13'b1111111111100, 13'b0000000000000, 13'b0000000000001, 13'b1111111111111, 13'b1111111111100, 13'b0000000000110, 13'b0000000001110, 13'b0000000001000, 13'b1111111110111, 13'b0000000000011, 13'b1111111111111, 13'b1111111111110, 13'b0000000000001, 13'b0000000000001, 13'b1111111111011, 13'b0000000000101, 13'b1111111111010, 13'b0000000000011, 13'b1111111111111, 13'b1111111101101, 13'b1111111111110, 13'b0000000001110}, 
{13'b1111111111110, 13'b1111111111010, 13'b0000000000100, 13'b0000000010000, 13'b0000000000101, 13'b0000000000101, 13'b0000000000010, 13'b1111111110011, 13'b1111111110010, 13'b0000000000100, 13'b0000000000000, 13'b0000000000010, 13'b0000000000001, 13'b0000000000000, 13'b0000000001101, 13'b0000000000000, 13'b1111111111100, 13'b0000000000110, 13'b1111111111110, 13'b1111111111101, 13'b0000000000111, 13'b1111111111000, 13'b1111111111110, 13'b0000000001000, 13'b0000000000001, 13'b1111111111001, 13'b1111111110011, 13'b1111111111111, 13'b1111111101110, 13'b0000000000011, 13'b0000000000110, 13'b0000000000000}, 
{13'b1111111111111, 13'b1111111111110, 13'b1111111111111, 13'b1111111111101, 13'b1111111110111, 13'b1111111110111, 13'b0000000000100, 13'b0000000000000, 13'b1111111110100, 13'b0000000001010, 13'b1111111111110, 13'b1111111111111, 13'b1111111111000, 13'b0000000000000, 13'b0000000000001, 13'b1111111111100, 13'b1111111111110, 13'b1111111111101, 13'b1111111111010, 13'b0000000000000, 13'b1111111110111, 13'b0000000000110, 13'b1111111110010, 13'b0000000000000, 13'b0000000000010, 13'b0000000000111, 13'b0000000000001, 13'b0000000000000, 13'b0000000010010, 13'b0000000000011, 13'b0000000000000, 13'b0000000000101}, 
{13'b1111111111110, 13'b0000000010000, 13'b1111111111111, 13'b1111111111101, 13'b1111111110010, 13'b1111111111011, 13'b0000000011010, 13'b1111111010011, 13'b1111111101001, 13'b1111111110011, 13'b1111111110001, 13'b1111111101111, 13'b1111111111111, 13'b0000000011110, 13'b1111111111110, 13'b0000000000000, 13'b1111111110010, 13'b0000000011100, 13'b1111111100101, 13'b0000000000000, 13'b1111111111111, 13'b1111111101010, 13'b0000000000000, 13'b1111111111111, 13'b0000000000011, 13'b1111111111100, 13'b1111111110110, 13'b1111111111111, 13'b0000000001011, 13'b0000000000000, 13'b1111111111010, 13'b0000000000000}, 
{13'b0000000010111, 13'b1111111111000, 13'b0000000001000, 13'b1111111111101, 13'b0000000000100, 13'b1111111111111, 13'b1111111111111, 13'b1111111111010, 13'b0000000000000, 13'b0000000000101, 13'b1111111111111, 13'b1111111111100, 13'b1111111111111, 13'b0000000001110, 13'b0000000000001, 13'b0000000000010, 13'b0000000000001, 13'b1111111111110, 13'b0000000000001, 13'b0000000000000, 13'b1111111111111, 13'b1111111111111, 13'b1111111101100, 13'b1111111111111, 13'b0000000000011, 13'b1111111111000, 13'b1111111110111, 13'b1111111111111, 13'b1111111111111, 13'b0000000100011, 13'b1111111101101, 13'b1111111111000}, 
{13'b1111111111101, 13'b1111111111001, 13'b1111111111011, 13'b0000000000010, 13'b0000000001000, 13'b1111111110111, 13'b1111111111111, 13'b1111111110001, 13'b0000000000011, 13'b0000000001000, 13'b1111111110010, 13'b1111111101111, 13'b0000000000001, 13'b1111111010100, 13'b1111111111011, 13'b1111111111000, 13'b1111111110011, 13'b1111111111111, 13'b0000000001000, 13'b0000000000000, 13'b1111111111101, 13'b1111111111101, 13'b0000000000000, 13'b0000000000000, 13'b1111111111100, 13'b1111111001111, 13'b1111111011100, 13'b1111111101110, 13'b0000000000011, 13'b0000000001101, 13'b1111111111111, 13'b0000000001111}, 
{13'b1111111111010, 13'b1111111110010, 13'b0000000001010, 13'b0000000000100, 13'b0000000000010, 13'b1111111111010, 13'b1111111111101, 13'b0000000000110, 13'b0000000100010, 13'b1111111110101, 13'b1111111111111, 13'b1111111111111, 13'b0000000000111, 13'b1111111111100, 13'b1111111111110, 13'b1111111111110, 13'b1111111111001, 13'b1111111111111, 13'b0000000000000, 13'b0000000001110, 13'b1111111110111, 13'b1111111111111, 13'b0000000001000, 13'b1111111111111, 13'b0000000000000, 13'b0000000100001, 13'b0000000010100, 13'b0000000000000, 13'b0000000000000, 13'b1111111100101, 13'b1111111111011, 13'b1111111111111}, 
{13'b0000000000000, 13'b0000000000011, 13'b1111111111111, 13'b0000000000000, 13'b0000000001110, 13'b1111111100001, 13'b0000000000000, 13'b1111111111001, 13'b0000000001011, 13'b0000000000000, 13'b1111111111110, 13'b0000000000000, 13'b0000000000000, 13'b1111111111111, 13'b0000000000000, 13'b1111111111001, 13'b0000000010000, 13'b1111111111111, 13'b1111111111111, 13'b1111111111111, 13'b0000000000000, 13'b1111111111111, 13'b0000000000000, 13'b1111111111111, 13'b0000000000000, 13'b1111111101011, 13'b0000000000011, 13'b0000000001011, 13'b1111111111111, 13'b0000000000110, 13'b1111111111111, 13'b0000000000100}, 
{13'b1111111110011, 13'b0000000000000, 13'b1111111100001, 13'b0000000000000, 13'b1111111111100, 13'b1111111111101, 13'b1111111111111, 13'b1111111111010, 13'b1111111111101, 13'b1111111111011, 13'b0000000000011, 13'b0000000000001, 13'b1111111110100, 13'b0000000000000, 13'b1111111111111, 13'b1111111111111, 13'b0000000000100, 13'b1111111111110, 13'b1111111111110, 13'b1111111111110, 13'b1111111111111, 13'b0000000010001, 13'b1111111111111, 13'b0000000000000, 13'b1111111111111, 13'b0000000010100, 13'b0000000001100, 13'b0000000000010, 13'b1111111111001, 13'b1111111111111, 13'b0000000000100, 13'b0000000000011}, 
{13'b0000000000010, 13'b0000000000010, 13'b1111111111111, 13'b0000000000000, 13'b1111111100010, 13'b0000000000010, 13'b0000000000001, 13'b1111111111111, 13'b0000000000000, 13'b1111111110101, 13'b1111111111111, 13'b0000000000000, 13'b1111111110101, 13'b0000000000000, 13'b0000000000000, 13'b0000000000000, 13'b0000000000000, 13'b1111111101001, 13'b0000000000000, 13'b1111111111111, 13'b1111111111111, 13'b0000000000000, 13'b0000000001000, 13'b1111111111111, 13'b0000000000000, 13'b0000000011101, 13'b0000000010101, 13'b0000000000000, 13'b0000000000000, 13'b1111111110001, 13'b0000000000000, 13'b1111111111111}, 
{13'b0000000000100, 13'b0000000000011, 13'b0000000010000, 13'b1111111110000, 13'b0000000001000, 13'b0000000000111, 13'b0000000000000, 13'b0000000001100, 13'b0000000000000, 13'b1111111111111, 13'b0000000000010, 13'b0000000000000, 13'b1111111111111, 13'b0000000000111, 13'b1111111111111, 13'b1111111111101, 13'b0000000000000, 13'b0000000000010, 13'b1111111111100, 13'b0000000000110, 13'b0000000000010, 13'b1111111011010, 13'b1111111111000, 13'b0000000000101, 13'b1111111111111, 13'b1111111011111, 13'b1111111110111, 13'b1111111111110, 13'b1111111111111, 13'b1111111111100, 13'b0000000000000, 13'b1111111111101}, 
{13'b0000000000000, 13'b1111111111111, 13'b1111111111010, 13'b1111111110101, 13'b0000000000010, 13'b0000000000000, 13'b0000000000110, 13'b1111111111111, 13'b0000000001111, 13'b1111111111111, 13'b0000000000000, 13'b1111111101010, 13'b1111111111111, 13'b0000000001000, 13'b1111111111111, 13'b1111111101111, 13'b0000000000000, 13'b1111111111111, 13'b0000000010000, 13'b1111111111111, 13'b1111111100100, 13'b1111111111111, 13'b0000000010000, 13'b1111111111111, 13'b1111111111111, 13'b0000000001000, 13'b1111111111001, 13'b0000000000100, 13'b0000000000000, 13'b1111111110011, 13'b0000000000000, 13'b0000000000000}, 
{13'b1111111110010, 13'b0000000000000, 13'b0000000000000, 13'b1111111111111, 13'b0000000011111, 13'b1111111111000, 13'b1111111111111, 13'b1111111111111, 13'b1111111111101, 13'b1111111111100, 13'b0000000000100, 13'b0000000001000, 13'b1111111111101, 13'b0000000001111, 13'b0000000000000, 13'b1111111111111, 13'b1111111101101, 13'b1111111111111, 13'b0000000000000, 13'b1111111111010, 13'b0000000000000, 13'b0000000000010, 13'b0000000000000, 13'b1111111111111, 13'b1111111111100, 13'b1111111110011, 13'b1111111101101, 13'b0000000000000, 13'b1111111111000, 13'b0000000000010, 13'b1111111111111, 13'b0000000000100}, 
{13'b1111111100101, 13'b1111111110101, 13'b1111111110110, 13'b0000000000000, 13'b0000000100100, 13'b1111111110001, 13'b0000000000000, 13'b1111111111100, 13'b1111111100101, 13'b0000000001000, 13'b1111111111111, 13'b0000000100100, 13'b0000000000000, 13'b1111111111100, 13'b1111111111111, 13'b0000000000010, 13'b1111111111110, 13'b0000000000000, 13'b1111111111101, 13'b0000000011111, 13'b0000000000010, 13'b1111111111101, 13'b0000000000111, 13'b1111111111111, 13'b1111111111111, 13'b1111111111001, 13'b1111111111101, 13'b1111111100010, 13'b1111111110110, 13'b1111111111111, 13'b1111111111111, 13'b1111111111100}, 
{13'b0000000001110, 13'b1111111001100, 13'b1111111010001, 13'b1111111110101, 13'b0000000101010, 13'b1111111111111, 13'b1111111101001, 13'b0000000010000, 13'b0000000000011, 13'b0000000000000, 13'b0000000001101, 13'b1111111101110, 13'b0000000000000, 13'b0000000000000, 13'b1111111111101, 13'b0000000000001, 13'b1111111111001, 13'b1111111000101, 13'b0000000001010, 13'b0000000010110, 13'b0000000010000, 13'b0000000000000, 13'b0000000000001, 13'b1111111100110, 13'b1111111010111, 13'b1111111111111, 13'b1111111101100, 13'b1111111100010, 13'b1111111110011, 13'b1111111000111, 13'b0000000011010, 13'b0000000011011}, 
{13'b0000000000000, 13'b0000000000000, 13'b0000000000000, 13'b0000000000000, 13'b0000000010000, 13'b1111111110100, 13'b0000000000001, 13'b0000000000100, 13'b1111111101001, 13'b0000000000010, 13'b1111111111111, 13'b1111111111111, 13'b1111111111111, 13'b0000000001111, 13'b0000000000011, 13'b0000000000001, 13'b0000000000011, 13'b0000000010101, 13'b1111111110010, 13'b0000000000000, 13'b1111111110101, 13'b1111111111111, 13'b0000000010100, 13'b0000000000000, 13'b1111111111111, 13'b1111111011100, 13'b1111111111111, 13'b1111111110110, 13'b1111111111100, 13'b0000000000000, 13'b0000000001000, 13'b0000000000110}, 
{13'b1111111111101, 13'b0000000001000, 13'b1111111101100, 13'b0000000000001, 13'b0000000001100, 13'b1111111111101, 13'b1111111111111, 13'b0000000001010, 13'b0000000000000, 13'b1111111111111, 13'b1111111111011, 13'b0000000000000, 13'b0000000000000, 13'b1111111111101, 13'b1111111111000, 13'b1111111111011, 13'b1111111111100, 13'b1111111111011, 13'b1111111111000, 13'b0000000000000, 13'b1111111111111, 13'b1111111111101, 13'b1111111111011, 13'b0000000011001, 13'b0000000000000, 13'b1111111101000, 13'b1111111111111, 13'b0000000000111, 13'b0000000000000, 13'b0000000000000, 13'b0000000010000, 13'b1111111111111}, 
{13'b1111111111111, 13'b0000000000000, 13'b1111111111111, 13'b1111111110110, 13'b1111111001000, 13'b0000000000000, 13'b0000000000000, 13'b1111111111111, 13'b1111111011001, 13'b0000000000101, 13'b1111111111001, 13'b1111111111111, 13'b0000000000000, 13'b1111111101000, 13'b1111111111101, 13'b1111111111111, 13'b0000000000000, 13'b0000000000000, 13'b0000000000010, 13'b0000000010110, 13'b1111111111000, 13'b1111111101100, 13'b0000000000000, 13'b1111111101111, 13'b1111111111001, 13'b1111111110001, 13'b1111111111111, 13'b1111111111111, 13'b1111111111110, 13'b1111111100001, 13'b1111111111101, 13'b0000000001111}, 
{13'b0000000000111, 13'b0000000001110, 13'b1111111111111, 13'b0000000001010, 13'b1111111110010, 13'b1111111111000, 13'b0000000000110, 13'b0000000000100, 13'b1111111111100, 13'b1111111111111, 13'b1111111111111, 13'b1111111111111, 13'b1111111111111, 13'b1111111101011, 13'b1111111111111, 13'b0000000001001, 13'b1111111111000, 13'b0000000000010, 13'b1111111111111, 13'b1111111111111, 13'b0000000001101, 13'b1111111101011, 13'b0000000010001, 13'b0000000000011, 13'b0000000000000, 13'b0000000001101, 13'b0000000000000, 13'b1111111111101, 13'b1111111100111, 13'b1111111111000, 13'b1111111110101, 13'b0000000001011}, 
{13'b0000000000000, 13'b0000000000000, 13'b1111111101000, 13'b1111111111111, 13'b0000000001101, 13'b1111111110110, 13'b1111111111111, 13'b1111111111111, 13'b0000000000001, 13'b0000000000000, 13'b0000000000000, 13'b1111111110010, 13'b0000000000110, 13'b0000000000000, 13'b0000000000000, 13'b0000000000010, 13'b1111111111111, 13'b1111111110110, 13'b0000000000001, 13'b0000000000000, 13'b1111111111101, 13'b1111111111110, 13'b0000000010010, 13'b1111111111111, 13'b0000000000000, 13'b1111111101101, 13'b1111111101011, 13'b0000000001111, 13'b1111111111111, 13'b1111111111111, 13'b0000000000001, 13'b0000000010010}, 
{13'b1111111101010, 13'b1111111111111, 13'b1111111110010, 13'b0000000000000, 13'b1111111101001, 13'b0000000000000, 13'b1111111111111, 13'b1111111111011, 13'b1111111011101, 13'b1111111111110, 13'b0000000000000, 13'b1111111111111, 13'b1111111111111, 13'b0000000000000, 13'b1111111111111, 13'b1111111111100, 13'b1111111110110, 13'b1111111111001, 13'b0000000000100, 13'b1111111111111, 13'b1111111111110, 13'b0000000000000, 13'b0000000010101, 13'b1111111111111, 13'b0000000001001, 13'b0000000000101, 13'b1111111110111, 13'b0000000001101, 13'b1111111111101, 13'b0000000000000, 13'b1111111111111, 13'b0000000100101}, 
{13'b1111111101011, 13'b0000000000001, 13'b0000000000011, 13'b1111111111110, 13'b0000000001111, 13'b1111111101100, 13'b1111111111111, 13'b0000000010000, 13'b0000000001010, 13'b0000000000000, 13'b1111111111111, 13'b1111111111011, 13'b1111111111010, 13'b1111111111011, 13'b1111111111100, 13'b0000000000101, 13'b1111111111111, 13'b0000000000000, 13'b0000000001001, 13'b0000000000000, 13'b0000000000000, 13'b0000000000000, 13'b0000000010000, 13'b0000000000010, 13'b0000000000000, 13'b1111111111001, 13'b1111111111111, 13'b0000000000000, 13'b1111111111111, 13'b1111111111111, 13'b1111111111111, 13'b0000000000100}, 
{13'b1111111111111, 13'b0000000000000, 13'b1111111110010, 13'b1111111111011, 13'b0000000010010, 13'b1111111111111, 13'b1111111111011, 13'b0000000001111, 13'b1111111111100, 13'b0000000010010, 13'b0000000000101, 13'b1111111111000, 13'b0000000000000, 13'b0000000000000, 13'b1111111111111, 13'b0000000000001, 13'b1111111111011, 13'b1111111101111, 13'b0000000010001, 13'b0000000001001, 13'b0000000101000, 13'b0000000001100, 13'b0000000001111, 13'b1111111111111, 13'b0000000000000, 13'b0000000000000, 13'b0000000000011, 13'b0000000000101, 13'b1111111100101, 13'b1111111111111, 13'b1111111111111, 13'b1111111111111}, 
{13'b0000000000000, 13'b1111111111010, 13'b1111111111001, 13'b0000000000000, 13'b1111111110000, 13'b0000000000000, 13'b0000000001100, 13'b0000000000110, 13'b0000000000011, 13'b1111111111001, 13'b0000000000000, 13'b1111111111111, 13'b1111111111111, 13'b1111111111111, 13'b1111111111101, 13'b0000000001100, 13'b1111111111111, 13'b1111111111111, 13'b1111111101100, 13'b0000000000000, 13'b1111111110011, 13'b1111111111111, 13'b0000000000000, 13'b1111111111111, 13'b0000000000000, 13'b0000000000001, 13'b0000000000001, 13'b0000000001000, 13'b1111111111011, 13'b1111111111111, 13'b1111111100011, 13'b0000000000101}, 
{13'b0000000011100, 13'b1111111111111, 13'b0000000000100, 13'b1111111111001, 13'b1111111111010, 13'b0000000000010, 13'b0000000001010, 13'b0000000000000, 13'b0000000100001, 13'b0000000000000, 13'b1111111111110, 13'b0000000000001, 13'b0000000000110, 13'b1111111111111, 13'b0000000000011, 13'b0000000000110, 13'b1111111111111, 13'b1111111100011, 13'b1111111111100, 13'b1111111111111, 13'b0000000000111, 13'b0000000000000, 13'b1111111111111, 13'b0000000000111, 13'b0000000000001, 13'b1111111101111, 13'b1111111111001, 13'b0000000001000, 13'b1111111111110, 13'b0000000010000, 13'b1111111111111, 13'b1111111110100}, 
{13'b0000000000000, 13'b0000000000110, 13'b1111111111111, 13'b1111111111101, 13'b1111111101001, 13'b1111111111111, 13'b0000000000010, 13'b1111111111101, 13'b0000000001010, 13'b1111111111101, 13'b1111111111111, 13'b1111111111101, 13'b1111111111111, 13'b1111111111101, 13'b0000000000000, 13'b0000000010100, 13'b0000000000000, 13'b1111111111111, 13'b1111111111111, 13'b1111111111111, 13'b1111111111111, 13'b1111111111111, 13'b0000000000010, 13'b0000000001000, 13'b0000000000000, 13'b0000000000000, 13'b0000000000010, 13'b1111111111111, 13'b0000000000000, 13'b0000000000001, 13'b0000000000000, 13'b0000000000110}, 
{13'b1111111101100, 13'b0000000001000, 13'b0000000000001, 13'b1111111111001, 13'b1111111100110, 13'b1111111111110, 13'b0000000000100, 13'b1111111100110, 13'b0000000100000, 13'b0000000000100, 13'b0000000000001, 13'b0000000000110, 13'b0000000000010, 13'b0000000000000, 13'b0000000011010, 13'b1111111111010, 13'b0000000000000, 13'b0000000000000, 13'b1111111111111, 13'b0000000000000, 13'b1111111100100, 13'b0000000000001, 13'b0000000001001, 13'b0000000000010, 13'b0000000000010, 13'b1111111010101, 13'b1111111101010, 13'b1111111110000, 13'b0000000000000, 13'b1111111111111, 13'b0000000010100, 13'b1111111110010}, 
{13'b1111111111111, 13'b1111111110011, 13'b1111111111001, 13'b1111111100101, 13'b1111111101111, 13'b0000000010101, 13'b0000000010011, 13'b1111111110101, 13'b0000000000010, 13'b1111111111101, 13'b1111111111001, 13'b1111111101111, 13'b0000000000110, 13'b1111111101101, 13'b0000000001100, 13'b1111111111111, 13'b0000000010101, 13'b1111111111111, 13'b1111111111111, 13'b1111111110111, 13'b1111111111101, 13'b1111111111011, 13'b1111111101110, 13'b0000000000101, 13'b1111111111111, 13'b1111111111111, 13'b1111111110001, 13'b0000000010100, 13'b0000000010001, 13'b1111111111010, 13'b1111111010111, 13'b0000000001001}, 
{13'b0000000000000, 13'b1111111111110, 13'b1111111111111, 13'b1111111111001, 13'b0000000000001, 13'b0000000000000, 13'b0000000000100, 13'b0000000000000, 13'b0000000000111, 13'b1111111111111, 13'b0000000000000, 13'b0000000000110, 13'b0000000000000, 13'b0000000000000, 13'b1111111110111, 13'b1111111111001, 13'b0000000000000, 13'b0000000001011, 13'b0000000000011, 13'b0000000001000, 13'b1111111111110, 13'b1111111110101, 13'b1111111111111, 13'b0000000000100, 13'b1111111111111, 13'b0000000000010, 13'b1111111111111, 13'b0000000000100, 13'b0000000000000, 13'b0000000000101, 13'b1111111100111, 13'b1111111111111}, 
{13'b0000000010011, 13'b1111111111111, 13'b0000000001001, 13'b1111111101100, 13'b1111111110011, 13'b1111111111111, 13'b1111111111111, 13'b0000000000001, 13'b0000000000000, 13'b1111111110111, 13'b0000000000000, 13'b0000000000000, 13'b0000000000000, 13'b0000000000000, 13'b1111111110111, 13'b0000000001001, 13'b1111111111111, 13'b1111111111110, 13'b0000000000000, 13'b0000000000111, 13'b1111111110011, 13'b0000000000111, 13'b0000000001000, 13'b0000000001000, 13'b1111111111111, 13'b0000000100011, 13'b1111111110110, 13'b0000000010111, 13'b1111111111100, 13'b1111111101000, 13'b1111111110100, 13'b0000000001000}, 
{13'b1111111011101, 13'b1111111111110, 13'b1111111110110, 13'b1111111111111, 13'b0000000010000, 13'b1111111110100, 13'b1111111111100, 13'b0000000001111, 13'b0000000000110, 13'b1111111110000, 13'b0000000000000, 13'b1111111111110, 13'b1111111111111, 13'b0000000001000, 13'b1111111110000, 13'b1111111111111, 13'b0000000000000, 13'b1111111111111, 13'b1111111111110, 13'b0000000000000, 13'b1111111110011, 13'b1111111111111, 13'b0000000000000, 13'b1111111101010, 13'b0000000000100, 13'b0000000100111, 13'b0000000010110, 13'b1111111111101, 13'b1111111110101, 13'b1111111100011, 13'b0000000000000, 13'b1111111111100}, 
{13'b0000000000001, 13'b0000000001101, 13'b0000000000001, 13'b1111111110110, 13'b0000000000000, 13'b1111111111110, 13'b0000000000000, 13'b0000000001101, 13'b0000000001101, 13'b1111111110111, 13'b0000000001000, 13'b0000000000001, 13'b1111111111111, 13'b1111111111111, 13'b1111111110101, 13'b0000000010000, 13'b1111111111101, 13'b1111111101011, 13'b0000000000111, 13'b1111111111111, 13'b1111111111111, 13'b0000000000111, 13'b1111111111011, 13'b1111111111111, 13'b1111111111100, 13'b0000000000101, 13'b1111111110111, 13'b0000000001000, 13'b1111111101000, 13'b0000000000101, 13'b1111111111111, 13'b0000000001010}, 
{13'b1111111111101, 13'b0000000000000, 13'b0000000000101, 13'b0000000000000, 13'b1111111111100, 13'b1111111111111, 13'b0000000000110, 13'b1111111111111, 13'b0000000000000, 13'b0000000000000, 13'b0000000000000, 13'b0000000000001, 13'b1111111111001, 13'b0000000000000, 13'b0000000000111, 13'b0000000000010, 13'b0000000000110, 13'b1111111111111, 13'b1111111111111, 13'b0000000001000, 13'b0000000001111, 13'b1111111111001, 13'b0000000000000, 13'b1111111111111, 13'b0000000000000, 13'b1111111100010, 13'b1111111111111, 13'b1111111111011, 13'b1111111111111, 13'b0000000100100, 13'b0000000000000, 13'b1111111110010}, 
{13'b1111111111110, 13'b1111111111000, 13'b1111111111111, 13'b0000000000000, 13'b0000000000101, 13'b1111111111111, 13'b0000000000000, 13'b1111111111110, 13'b0000000000100, 13'b1111111111111, 13'b0000000000000, 13'b0000000000010, 13'b0000000010010, 13'b1111111111001, 13'b0000000000000, 13'b1111111001001, 13'b1111111111111, 13'b1111111111100, 13'b0000000000000, 13'b1111111111100, 13'b0000000000101, 13'b1111111110001, 13'b0000000000111, 13'b0000000000110, 13'b1111111111111, 13'b1111111010010, 13'b1111111110001, 13'b1111111111110, 13'b1111111111110, 13'b0000000011000, 13'b1111111111111, 13'b0000000001001}, 
{13'b0000000000011, 13'b0000000000000, 13'b0000000001011, 13'b1111111111000, 13'b1111111111011, 13'b0000000001111, 13'b1111111110101, 13'b0000000000011, 13'b1111111101100, 13'b0000000000000, 13'b0000000000001, 13'b1111111111010, 13'b0000000000000, 13'b0000000000000, 13'b1111111110011, 13'b0000000011011, 13'b1111111110000, 13'b1111111111111, 13'b0000000000111, 13'b1111111111111, 13'b0000000000100, 13'b1111111100001, 13'b0000000010100, 13'b1111111111111, 13'b1111111111000, 13'b0000000011111, 13'b0000000001001, 13'b1111111110101, 13'b1111111110111, 13'b1111111011101, 13'b1111111111111, 13'b0000000000001}, 
{13'b1111111111111, 13'b0000000000000, 13'b1111111111101, 13'b1111111101110, 13'b1111111111111, 13'b1111111100110, 13'b0000000000000, 13'b0000000010011, 13'b0000000001111, 13'b0000000000001, 13'b0000000000000, 13'b1111111111000, 13'b0000000010101, 13'b1111111111111, 13'b1111111111111, 13'b1111111111111, 13'b0000000011011, 13'b0000000000000, 13'b1111111111101, 13'b1111111111100, 13'b1111111101011, 13'b0000000001000, 13'b0000000000000, 13'b0000000000000, 13'b0000000000010, 13'b1111111111011, 13'b1111111100010, 13'b0000000010001, 13'b1111111100011, 13'b0000000000011, 13'b1111111111010, 13'b0000000000000}, 
{13'b0000000000011, 13'b0000000001011, 13'b0000000000000, 13'b1111111111111, 13'b1111111100010, 13'b0000000000000, 13'b1111111111111, 13'b0000000001111, 13'b0000000010001, 13'b1111111111111, 13'b1111111111111, 13'b1111111111111, 13'b0000000000000, 13'b0000000000000, 13'b0000000000000, 13'b0000000000000, 13'b0000000000000, 13'b1111111111111, 13'b0000000001010, 13'b1111111111001, 13'b1111111100100, 13'b1111111111101, 13'b1111111111001, 13'b1111111111001, 13'b1111111111011, 13'b1111111111111, 13'b1111111111011, 13'b1111111111110, 13'b1111111111111, 13'b0000000001001, 13'b1111111111111, 13'b0000000011101}
};

localparam logic signed [12:0] bias [32] = '{
13'b0000001011110,  // 1.474280834197998
13'b0000000101100,  // 0.6914801001548767
13'b0000001011100,  // 1.4406442642211914
13'b0000001011010,  // 1.408045768737793
13'b0000000111111,  // 0.9864811301231384
13'b0000000110111,  // 0.8636202812194824
13'b1111111011000,  // -0.6153604388237
13'b0000000011110,  // 0.4839226007461548
13'b0000000011111,  // 0.4862793982028961
13'b0000000010111,  // 0.37162142992019653
13'b0000000011101,  // 0.45989668369293213
13'b0000001010011,  // 1.2998151779174805
13'b1111110111110,  // -1.016528844833374
13'b1111111101001,  // -0.35249894857406616
13'b0000000011100,  // 0.44582197070121765
13'b1111111111000,  // -0.1119980737566948
13'b1111111111011,  // -0.06717441976070404
13'b0000000000000,  // 0.00487547367811203
13'b0000000001100,  // 0.1946917623281479
13'b1111111001110,  // -0.7796769738197327
13'b0000000101110,  // 0.7287401556968689
13'b0000001101101,  // 1.714877724647522
13'b1111110011001,  // -1.5971007347106934
13'b0000000000100,  // 0.07393483817577362
13'b0000000010100,  // 0.3225609362125397
13'b0000000110110,  // 0.8453295230865479
13'b0000000111001,  // 0.898597240447998
13'b0000000010000,  // 0.2548799514770508
13'b0000000111110,  // 0.9735668301582336
13'b0000001001000,  // 1.1261906623840332
13'b0000000011100,  // 0.44768181443214417
13'b1111101101000   // -2.3676068782806396
};
endpackage