// Width: 11
// NFRAC: 5
package dense_2_11_5;

localparam logic signed [10:0] weights [64][32] = '{ 
{11'b00000001000, 11'b00000000000, 11'b11111111001, 11'b11111111111, 11'b00000001000, 11'b00000000000, 11'b11111111011, 11'b11111111111, 11'b11111110111, 11'b00000000010, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b11111111001, 11'b11111111110, 11'b11111110111, 11'b00000000000, 11'b11111111111, 11'b11111111001, 11'b11111111010, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b00000000011, 11'b00000001100, 11'b00000000101, 11'b11111111111, 11'b00000000001, 11'b11111110010, 11'b00000000000}, 
{11'b11111111100, 11'b11111111011, 11'b11111111011, 11'b11111111110, 11'b11111111111, 11'b00000000001, 11'b11111111000, 11'b00000000000, 11'b00000000000, 11'b11111111101, 11'b00000000100, 11'b11111111110, 11'b11111111110, 11'b11111111001, 11'b00000000000, 11'b11111111110, 11'b00000000000, 11'b11111111001, 11'b00000000101, 11'b00000000111, 11'b11111111110, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b11111111101, 11'b00000001000, 11'b00000000111, 11'b00000000000, 11'b00000000000, 11'b11111110000, 11'b00000000000, 11'b00000000000}, 
{11'b00000000010, 11'b11111111100, 11'b11111111011, 11'b11111111110, 11'b11111111101, 11'b11111111101, 11'b11111111010, 11'b00000000000, 11'b11111111011, 11'b00000000000, 11'b00000000000, 11'b11111111101, 11'b00000000010, 11'b11111111101, 11'b11111111111, 11'b11111111110, 11'b00000000000, 11'b00000000011, 11'b00000000001, 11'b00000000111, 11'b00000000001, 11'b11111111101, 11'b00000000000, 11'b00000000001, 11'b11111111111, 11'b00000000110, 11'b00000000100, 11'b00000000011, 11'b11111111111, 11'b11111111011, 11'b11111111111, 11'b00000000011}, 
{11'b00000000100, 11'b00000000000, 11'b00000000001, 11'b11111111111, 11'b11111101111, 11'b00000000000, 11'b00000000000, 11'b00000000111, 11'b00000000111, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b00000000110, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b11111111010, 11'b11111111110, 11'b00000000001, 11'b11111111101, 11'b11111111111, 11'b00000000000, 11'b11111111110, 11'b00000000010, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b11111111001, 11'b00000001001}, 
{11'b11111101010, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b11111111110, 11'b11111111011, 11'b00000000001, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b00000000110, 11'b00000000000, 11'b00000001010, 11'b11111111111, 11'b00000000110, 11'b11111110011, 11'b00000000000, 11'b11111111100, 11'b00000000101, 11'b00000001000, 11'b00000000000, 11'b00000000001, 11'b00000000101, 11'b00000000111, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b00000000111}, 
{11'b00000000001, 11'b11111111111, 11'b00000000100, 11'b11111101011, 11'b11111010011, 11'b11111110100, 11'b00000001011, 11'b11111101100, 11'b11111111111, 11'b11111101010, 11'b11111101111, 11'b11111110101, 11'b00000001011, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b11111111011, 11'b11111111111, 11'b11111110000, 11'b00000000000, 11'b00000000101, 11'b11111111111, 11'b00000000000, 11'b00000001000, 11'b00000000001, 11'b11111111111, 11'b11111111111, 11'b00000000110, 11'b11111111110, 11'b00000000110}, 
{11'b11111111110, 11'b11111111010, 11'b11111111000, 11'b11111111110, 11'b11111110110, 11'b00000000010, 11'b11111111010, 11'b11111111011, 11'b11111110010, 11'b00000000001, 11'b11111111111, 11'b11111111010, 11'b00000000011, 11'b11111111111, 11'b11111111110, 11'b11111101110, 11'b11111111111, 11'b00000000010, 11'b00000000110, 11'b11111111010, 11'b11111111011, 11'b11111111101, 11'b11111111111, 11'b00000000000, 11'b11111111110, 11'b11111101011, 11'b11111110111, 11'b11111111110, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b11111111111}, 
{11'b11111111011, 11'b11111111101, 11'b11111111101, 11'b11111111000, 11'b11111111100, 11'b11111111111, 11'b00000000011, 11'b11111111101, 11'b00000000110, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b00000000111, 11'b00000000000, 11'b11111111111, 11'b11111111101, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b00000000001, 11'b11111111010, 11'b00000000000, 11'b11111111111, 11'b11111111101, 11'b11111111111, 11'b00000000000, 11'b11111111111}, 
{11'b11111110000, 11'b11111111110, 11'b11111110011, 11'b00000000011, 11'b00000001111, 11'b11111111111, 11'b11111111111, 11'b00000000111, 11'b11111110001, 11'b11111111110, 11'b00000000000, 11'b11111111001, 11'b11111111111, 11'b00000000010, 11'b11111111001, 11'b00000011000, 11'b11111111111, 11'b00000000001, 11'b00000000110, 11'b00000000111, 11'b00000000000, 11'b11111110101, 11'b00000000000, 11'b00000001101, 11'b11111111010, 11'b00000010110, 11'b11111111011, 11'b11111111001, 11'b11111110000, 11'b11111110001, 11'b00000000000, 11'b00000000001}, 
{11'b00000000000, 11'b11111111111, 11'b11111111101, 11'b00000000000, 11'b00000001001, 11'b11111111111, 11'b11111111101, 11'b00000000010, 11'b00000000011, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b11111111100, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b00000000010, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b00000000001, 11'b11111111011, 11'b00000000010, 11'b00000000111, 11'b11111111111, 11'b00000000000, 11'b00000000001, 11'b00000000010}, 
{11'b00000000011, 11'b00000000000, 11'b11111111100, 11'b11111110111, 11'b11111100110, 11'b00000000100, 11'b00000000000, 11'b11111100101, 11'b00000000001, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b11111110011, 11'b11111111111, 11'b00000000111, 11'b00000000100, 11'b00000000110, 11'b11111110001, 11'b11111110100, 11'b00000000011, 11'b11111111110, 11'b11111111110, 11'b00000001011, 11'b11111111100, 11'b11111111111, 11'b11111111111, 11'b00000000110, 11'b11111111111, 11'b00000000000}, 
{11'b11111111001, 11'b11111110000, 11'b00000000000, 11'b11111111111, 11'b00000001010, 11'b11111110111, 11'b11111111000, 11'b00000000011, 11'b11111111111, 11'b00000000100, 11'b00000000010, 11'b11111111101, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b11111110111, 11'b00000000101, 11'b00000000000, 11'b00000001001, 11'b00000000010, 11'b00000000000, 11'b11111111110, 11'b00000000100, 11'b11111111101, 11'b11111110110, 11'b11111111111, 11'b00000000101, 11'b11111111111, 11'b00000000000, 11'b11111111100, 11'b00000000100, 11'b00000001000}, 
{11'b00000000000, 11'b00000000000, 11'b00000000111, 11'b00000000000, 11'b11111111110, 11'b00000000101, 11'b00000000010, 11'b11111111111, 11'b00000000000, 11'b11111111011, 11'b11111111110, 11'b11111111010, 11'b11111111111, 11'b00000000001, 11'b11111111101, 11'b00000011010, 11'b00000000000, 11'b11111111100, 11'b11111111001, 11'b11111111111, 11'b00000000110, 11'b00000000100, 11'b00000000000, 11'b11111111111, 11'b00000000111, 11'b00000001000, 11'b00000001111, 11'b00000000000, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b11111111101}, 
{11'b11111111011, 11'b00000000001, 11'b00000000001, 11'b11111111000, 11'b11111110111, 11'b00000001111, 11'b00000000001, 11'b00000000000, 11'b11111111010, 11'b11111111101, 11'b00000000100, 11'b00000000010, 11'b00000000000, 11'b11111111101, 11'b00000001001, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b11111111110, 11'b00000000010, 11'b00000000000, 11'b00000000011, 11'b11111111111, 11'b00000000000, 11'b00000010101, 11'b11111111110, 11'b11111111111, 11'b11111111111, 11'b11111111100, 11'b11111111110, 11'b00000000101}, 
{11'b00000000001, 11'b00000000010, 11'b00000001010, 11'b11111111110, 11'b00000000011, 11'b00000001011, 11'b00000000000, 11'b11111111111, 11'b00000000011, 11'b11111111100, 11'b11111111111, 11'b11111111100, 11'b00000000000, 11'b00000001100, 11'b11111111111, 11'b00000000000, 11'b00000000111, 11'b00000000000, 11'b00000000000, 11'b11111110101, 11'b11111111000, 11'b11111111110, 11'b11111111111, 11'b11111111011, 11'b11111111110, 11'b11111111101, 11'b11111111001, 11'b11111111001, 11'b00000000000, 11'b00000000011, 11'b11111110011, 11'b00000000000}, 
{11'b11111110110, 11'b00000000000, 11'b11111111111, 11'b11111111110, 11'b11111111111, 11'b00000000100, 11'b11111111101, 11'b00000001000, 11'b11111110100, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b11111111101, 11'b00000000010, 11'b00000000101, 11'b11111111111, 11'b11111110111, 11'b11111111110, 11'b00000000011, 11'b00000000010, 11'b00000000000, 11'b00000000000, 11'b00000000010, 11'b11111111000, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b11111111011}, 
{11'b11111110101, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b00000000011, 11'b00000000000, 11'b00000000001, 11'b00000000001, 11'b00000000010, 11'b00000000010, 11'b00000000101, 11'b00000000000, 11'b11111111100, 11'b00000000000, 11'b00000001100, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b00000000011, 11'b00000000100, 11'b00000000000, 11'b00000000001, 11'b11111111111, 11'b11111111110, 11'b00000000000, 11'b11111111101, 11'b11111111011, 11'b00000000110, 11'b11111111111, 11'b00000000001, 11'b11111111001}, 
{11'b00000000000, 11'b11111111111, 11'b00000000001, 11'b00000000000, 11'b00000011101, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b00000000011, 11'b11111111101, 11'b00000000000, 11'b00000000000, 11'b00000000000, 11'b00000000100, 11'b00000000000, 11'b11111111011, 11'b11111111111, 11'b11111111101, 11'b00000001010, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b00000000010, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b00000000001}, 
{11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b00000000001, 11'b11111111110, 11'b11111111100, 11'b11111111110, 11'b00000001000, 11'b00000000000, 11'b00000000011, 11'b11111111111, 11'b00000000010, 11'b11111111110, 11'b11111111010, 11'b11111111001, 11'b00000000000, 11'b11111111111, 11'b11111111110, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b00000000010, 11'b00000000001, 11'b11111111011, 11'b00000000011, 11'b11111111010, 11'b00000000000, 11'b00000000000, 11'b11111111010, 11'b00000000000, 11'b00000000001, 11'b11111111111}, 
{11'b11111111111, 11'b11111111100, 11'b00000000000, 11'b11111111110, 11'b00000000110, 11'b11111111111, 11'b11111111111, 11'b00000000011, 11'b11111110011, 11'b00000000000, 11'b11111111110, 11'b11111111111, 11'b00000001011, 11'b00000000111, 11'b11111111100, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b11111111011, 11'b11111111100, 11'b00000000100, 11'b00000000000, 11'b11111111011, 11'b00000000000, 11'b11111111101, 11'b11111111110, 11'b00000000100, 11'b00000000000, 11'b11111111000}, 
{11'b00000010100, 11'b00000001010, 11'b11111111000, 11'b00000000000, 11'b11111110100, 11'b00000000000, 11'b00000000111, 11'b00000000000, 11'b00000000111, 11'b11111111111, 11'b11111111011, 11'b11111111101, 11'b00000000100, 11'b00000000000, 11'b11111111100, 11'b00000000100, 11'b00000010001, 11'b11111111011, 11'b11111110110, 11'b00000000000, 11'b11111111111, 11'b11111111010, 11'b11111111111, 11'b11111111111, 11'b00000000010, 11'b11111110100, 11'b00000000010, 11'b11111111111, 11'b00000000000, 11'b00000000011, 11'b11111111111, 11'b00000000001}, 
{11'b11111111101, 11'b11111111001, 11'b11111111110, 11'b11111111010, 11'b11111111111, 11'b00000000001, 11'b00000000000, 11'b11111111111, 11'b00000000001, 11'b11111111111, 11'b00000000000, 11'b11111111001, 11'b00000000011, 11'b00000000010, 11'b11111111100, 11'b00000001110, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b00000001010, 11'b11111110000, 11'b11111111100, 11'b11111111110, 11'b11111111111, 11'b00000000110, 11'b11111111110, 11'b00000000000, 11'b00000001111, 11'b11111101111, 11'b11111110100, 11'b00000000000}, 
{11'b00000000000, 11'b11111111110, 11'b11111111111, 11'b00000000000, 11'b11111101000, 11'b11111101100, 11'b00000000000, 11'b11111111111, 11'b11111110111, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b11111111110, 11'b11111111110, 11'b11111111101, 11'b11111111011, 11'b00000001001, 11'b00000000000, 11'b00000000001, 11'b11111111111, 11'b11111111101, 11'b00000000000, 11'b11111111101, 11'b00000000111, 11'b11111101100, 11'b00000000111, 11'b11111111111, 11'b11111111111, 11'b00000000110, 11'b11111111111, 11'b00000000111}, 
{11'b11111111111, 11'b00000000000, 11'b11111111110, 11'b00000000010, 11'b00000000001, 11'b11111110101, 11'b00000000000, 11'b00000000010, 11'b00000010010, 11'b11111111111, 11'b00000000000, 11'b00000000001, 11'b00000001011, 11'b11111111110, 11'b00000000000, 11'b00000000011, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b11111110111, 11'b00000000001, 11'b00000000010, 11'b00000000000, 11'b11111111111, 11'b00000000110, 11'b00000000000, 11'b00000000100, 11'b11111110010, 11'b00000000011, 11'b00000001100, 11'b00000000000}, 
{11'b11111110100, 11'b00000000110, 11'b11111110111, 11'b00000000011, 11'b11111111100, 11'b00000000000, 11'b00000001111, 11'b11111111000, 11'b11111110110, 11'b00000000101, 11'b11111111000, 11'b11111111111, 11'b11111111111, 11'b00000001011, 11'b11111111111, 11'b11111110110, 11'b11111111111, 11'b00000001110, 11'b11111110000, 11'b11111111111, 11'b00000001010, 11'b11111110100, 11'b00000000001, 11'b11111111111, 11'b00000001000, 11'b11111101111, 11'b11111110100, 11'b11111111001, 11'b11111111111, 11'b00000000011, 11'b00000000000, 11'b00000000101}, 
{11'b11111111101, 11'b00000000001, 11'b11111111111, 11'b00000000100, 11'b11111111110, 11'b00000000111, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b00000010000, 11'b00000000000, 11'b00000000110, 11'b00000000000, 11'b11111111001, 11'b11111111101, 11'b11111111111, 11'b11111111111, 11'b00000000001, 11'b11111111111, 11'b11111111010, 11'b11111111111, 11'b00000001001, 11'b00000001001, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b11111111100}, 
{11'b11111111101, 11'b00000000000, 11'b00000001000, 11'b00000000000, 11'b00000000000, 11'b11111111100, 11'b00000000000, 11'b11111100100, 11'b00000000110, 11'b00000000000, 11'b00000000000, 11'b11111110100, 11'b00000000000, 11'b11111111011, 11'b11111111110, 11'b00000000000, 11'b00000000000, 11'b00000000000, 11'b00000000011, 11'b00000000000, 11'b11111111111, 11'b00000001010, 11'b00000001100, 11'b11111111000, 11'b11111111011, 11'b00000000111, 11'b11111110110, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b00000000101}, 
{11'b11111111100, 11'b11111111111, 11'b11111111000, 11'b11111111001, 11'b11111111111, 11'b11111111011, 11'b00000000000, 11'b00000000010, 11'b11111111000, 11'b11111111101, 11'b11111111110, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b11111111110, 11'b00000000011, 11'b00000000111, 11'b00000000100, 11'b11111111011, 11'b00000000001, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b11111111101, 11'b00000000010, 11'b11111111101, 11'b00000000001, 11'b11111111111, 11'b11111110110, 11'b11111111111, 11'b00000000111}, 
{11'b11111111111, 11'b11111111101, 11'b00000000010, 11'b00000001000, 11'b00000000010, 11'b00000000010, 11'b00000000001, 11'b11111111001, 11'b11111111001, 11'b00000000010, 11'b00000000000, 11'b00000000001, 11'b00000000000, 11'b00000000000, 11'b00000000110, 11'b00000000000, 11'b11111111110, 11'b00000000011, 11'b11111111111, 11'b11111111110, 11'b00000000011, 11'b11111111100, 11'b11111111111, 11'b00000000100, 11'b00000000000, 11'b11111111100, 11'b11111111001, 11'b11111111111, 11'b11111110111, 11'b00000000001, 11'b00000000011, 11'b00000000000}, 
{11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b11111111110, 11'b11111111011, 11'b11111111011, 11'b00000000010, 11'b00000000000, 11'b11111111010, 11'b00000000101, 11'b11111111111, 11'b11111111111, 11'b11111111100, 11'b00000000000, 11'b00000000000, 11'b11111111110, 11'b11111111111, 11'b11111111110, 11'b11111111101, 11'b00000000000, 11'b11111111011, 11'b00000000011, 11'b11111111001, 11'b00000000000, 11'b00000000001, 11'b00000000011, 11'b00000000000, 11'b00000000000, 11'b00000001001, 11'b00000000001, 11'b00000000000, 11'b00000000010}, 
{11'b11111111111, 11'b00000001000, 11'b11111111111, 11'b11111111110, 11'b11111111001, 11'b11111111101, 11'b00000001101, 11'b11111101001, 11'b11111110100, 11'b11111111001, 11'b11111111000, 11'b11111110111, 11'b11111111111, 11'b00000001111, 11'b11111111111, 11'b00000000000, 11'b11111111001, 11'b00000001110, 11'b11111110010, 11'b00000000000, 11'b11111111111, 11'b11111110101, 11'b00000000000, 11'b11111111111, 11'b00000000001, 11'b11111111110, 11'b11111111011, 11'b11111111111, 11'b00000000101, 11'b00000000000, 11'b11111111101, 11'b00000000000}, 
{11'b00000001011, 11'b11111111100, 11'b00000000100, 11'b11111111110, 11'b00000000010, 11'b11111111111, 11'b11111111111, 11'b11111111101, 11'b00000000000, 11'b00000000010, 11'b11111111111, 11'b11111111110, 11'b11111111111, 11'b00000000111, 11'b00000000000, 11'b00000000001, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b11111110110, 11'b11111111111, 11'b00000000001, 11'b11111111100, 11'b11111111011, 11'b11111111111, 11'b11111111111, 11'b00000010001, 11'b11111110110, 11'b11111111100}, 
{11'b11111111110, 11'b11111111100, 11'b11111111101, 11'b00000000001, 11'b00000000100, 11'b11111111011, 11'b11111111111, 11'b11111111000, 11'b00000000001, 11'b00000000100, 11'b11111111001, 11'b11111110111, 11'b00000000000, 11'b11111101010, 11'b11111111101, 11'b11111111100, 11'b11111111001, 11'b11111111111, 11'b00000000100, 11'b00000000000, 11'b11111111110, 11'b11111111110, 11'b00000000000, 11'b00000000000, 11'b11111111110, 11'b11111100111, 11'b11111101110, 11'b11111110111, 11'b00000000001, 11'b00000000110, 11'b11111111111, 11'b00000000111}, 
{11'b11111111101, 11'b11111111001, 11'b00000000101, 11'b00000000010, 11'b00000000001, 11'b11111111101, 11'b11111111110, 11'b00000000011, 11'b00000010001, 11'b11111111010, 11'b11111111111, 11'b11111111111, 11'b00000000011, 11'b11111111110, 11'b11111111111, 11'b11111111111, 11'b11111111100, 11'b11111111111, 11'b00000000000, 11'b00000000111, 11'b11111111011, 11'b11111111111, 11'b00000000100, 11'b11111111111, 11'b00000000000, 11'b00000010000, 11'b00000001010, 11'b00000000000, 11'b00000000000, 11'b11111110010, 11'b11111111101, 11'b11111111111}, 
{11'b00000000000, 11'b00000000001, 11'b11111111111, 11'b00000000000, 11'b00000000111, 11'b11111110000, 11'b00000000000, 11'b11111111100, 11'b00000000101, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b11111111100, 11'b00000001000, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b11111110101, 11'b00000000001, 11'b00000000101, 11'b11111111111, 11'b00000000011, 11'b11111111111, 11'b00000000010}, 
{11'b11111111001, 11'b00000000000, 11'b11111110000, 11'b00000000000, 11'b11111111110, 11'b11111111110, 11'b11111111111, 11'b11111111101, 11'b11111111110, 11'b11111111101, 11'b00000000001, 11'b00000000000, 11'b11111111010, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b00000000010, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b00000001000, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b00000001010, 11'b00000000110, 11'b00000000001, 11'b11111111100, 11'b11111111111, 11'b00000000010, 11'b00000000001}, 
{11'b00000000001, 11'b00000000001, 11'b11111111111, 11'b00000000000, 11'b11111110001, 11'b00000000001, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b11111111010, 11'b11111111111, 11'b00000000000, 11'b11111111010, 11'b00000000000, 11'b00000000000, 11'b00000000000, 11'b00000000000, 11'b11111110100, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b00000000100, 11'b11111111111, 11'b00000000000, 11'b00000001110, 11'b00000001010, 11'b00000000000, 11'b00000000000, 11'b11111111000, 11'b00000000000, 11'b11111111111}, 
{11'b00000000010, 11'b00000000001, 11'b00000001000, 11'b11111111000, 11'b00000000100, 11'b00000000011, 11'b00000000000, 11'b00000000110, 11'b00000000000, 11'b11111111111, 11'b00000000001, 11'b00000000000, 11'b11111111111, 11'b00000000011, 11'b11111111111, 11'b11111111110, 11'b00000000000, 11'b00000000001, 11'b11111111110, 11'b00000000011, 11'b00000000001, 11'b11111101101, 11'b11111111100, 11'b00000000010, 11'b11111111111, 11'b11111101111, 11'b11111111011, 11'b11111111111, 11'b11111111111, 11'b11111111110, 11'b00000000000, 11'b11111111110}, 
{11'b00000000000, 11'b11111111111, 11'b11111111101, 11'b11111111010, 11'b00000000001, 11'b00000000000, 11'b00000000011, 11'b11111111111, 11'b00000000111, 11'b11111111111, 11'b00000000000, 11'b11111110101, 11'b11111111111, 11'b00000000100, 11'b11111111111, 11'b11111110111, 11'b00000000000, 11'b11111111111, 11'b00000001000, 11'b11111111111, 11'b11111110010, 11'b11111111111, 11'b00000001000, 11'b11111111111, 11'b11111111111, 11'b00000000100, 11'b11111111100, 11'b00000000010, 11'b00000000000, 11'b11111111001, 11'b00000000000, 11'b00000000000}, 
{11'b11111111001, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b00000001111, 11'b11111111100, 11'b11111111111, 11'b11111111111, 11'b11111111110, 11'b11111111110, 11'b00000000010, 11'b00000000100, 11'b11111111110, 11'b00000000111, 11'b00000000000, 11'b11111111111, 11'b11111110110, 11'b11111111111, 11'b00000000000, 11'b11111111101, 11'b00000000000, 11'b00000000001, 11'b00000000000, 11'b11111111111, 11'b11111111110, 11'b11111111001, 11'b11111110110, 11'b00000000000, 11'b11111111100, 11'b00000000001, 11'b11111111111, 11'b00000000010}, 
{11'b11111110010, 11'b11111111010, 11'b11111111011, 11'b00000000000, 11'b00000010010, 11'b11111111000, 11'b00000000000, 11'b11111111110, 11'b11111110010, 11'b00000000100, 11'b11111111111, 11'b00000010010, 11'b00000000000, 11'b11111111110, 11'b11111111111, 11'b00000000001, 11'b11111111111, 11'b00000000000, 11'b11111111110, 11'b00000001111, 11'b00000000001, 11'b11111111110, 11'b00000000011, 11'b11111111111, 11'b11111111111, 11'b11111111100, 11'b11111111110, 11'b11111110001, 11'b11111111011, 11'b11111111111, 11'b11111111111, 11'b11111111110}, 
{11'b00000000111, 11'b11111100110, 11'b11111101000, 11'b11111111010, 11'b00000010101, 11'b11111111111, 11'b11111110100, 11'b00000001000, 11'b00000000001, 11'b00000000000, 11'b00000000110, 11'b11111110111, 11'b00000000000, 11'b00000000000, 11'b11111111110, 11'b00000000000, 11'b11111111100, 11'b11111100010, 11'b00000000101, 11'b00000001011, 11'b00000001000, 11'b00000000000, 11'b00000000000, 11'b11111110011, 11'b11111101011, 11'b11111111111, 11'b11111110110, 11'b11111110001, 11'b11111111001, 11'b11111100011, 11'b00000001101, 11'b00000001101}, 
{11'b00000000000, 11'b00000000000, 11'b00000000000, 11'b00000000000, 11'b00000001000, 11'b11111111010, 11'b00000000000, 11'b00000000010, 11'b11111110100, 11'b00000000001, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b00000000111, 11'b00000000001, 11'b00000000000, 11'b00000000001, 11'b00000001010, 11'b11111111001, 11'b00000000000, 11'b11111111010, 11'b11111111111, 11'b00000001010, 11'b00000000000, 11'b11111111111, 11'b11111101110, 11'b11111111111, 11'b11111111011, 11'b11111111110, 11'b00000000000, 11'b00000000100, 11'b00000000011}, 
{11'b11111111110, 11'b00000000100, 11'b11111110110, 11'b00000000000, 11'b00000000110, 11'b11111111110, 11'b11111111111, 11'b00000000101, 11'b00000000000, 11'b11111111111, 11'b11111111101, 11'b00000000000, 11'b00000000000, 11'b11111111110, 11'b11111111100, 11'b11111111101, 11'b11111111110, 11'b11111111101, 11'b11111111100, 11'b00000000000, 11'b11111111111, 11'b11111111110, 11'b11111111101, 11'b00000001100, 11'b00000000000, 11'b11111110100, 11'b11111111111, 11'b00000000011, 11'b00000000000, 11'b00000000000, 11'b00000001000, 11'b11111111111}, 
{11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b11111111011, 11'b11111100100, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b11111101100, 11'b00000000010, 11'b11111111100, 11'b11111111111, 11'b00000000000, 11'b11111110100, 11'b11111111110, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b00000000001, 11'b00000001011, 11'b11111111100, 11'b11111110110, 11'b00000000000, 11'b11111110111, 11'b11111111100, 11'b11111111000, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b11111110000, 11'b11111111110, 11'b00000000111}, 
{11'b00000000011, 11'b00000000111, 11'b11111111111, 11'b00000000101, 11'b11111111001, 11'b11111111100, 11'b00000000011, 11'b00000000010, 11'b11111111110, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b11111110101, 11'b11111111111, 11'b00000000100, 11'b11111111100, 11'b00000000001, 11'b11111111111, 11'b11111111111, 11'b00000000110, 11'b11111110101, 11'b00000001000, 11'b00000000001, 11'b00000000000, 11'b00000000110, 11'b00000000000, 11'b11111111110, 11'b11111110011, 11'b11111111100, 11'b11111111010, 11'b00000000101}, 
{11'b00000000000, 11'b00000000000, 11'b11111110100, 11'b11111111111, 11'b00000000110, 11'b11111111011, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b00000000000, 11'b11111111001, 11'b00000000011, 11'b00000000000, 11'b00000000000, 11'b00000000001, 11'b11111111111, 11'b11111111011, 11'b00000000000, 11'b00000000000, 11'b11111111110, 11'b11111111111, 11'b00000001001, 11'b11111111111, 11'b00000000000, 11'b11111110110, 11'b11111110101, 11'b00000000111, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b00000001001}, 
{11'b11111110101, 11'b11111111111, 11'b11111111001, 11'b00000000000, 11'b11111110100, 11'b00000000000, 11'b11111111111, 11'b11111111101, 11'b11111101110, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b11111111110, 11'b11111111011, 11'b11111111100, 11'b00000000010, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b00000001010, 11'b11111111111, 11'b00000000100, 11'b00000000010, 11'b11111111011, 11'b00000000110, 11'b11111111110, 11'b00000000000, 11'b11111111111, 11'b00000010010}, 
{11'b11111110101, 11'b00000000000, 11'b00000000001, 11'b11111111111, 11'b00000000111, 11'b11111110110, 11'b11111111111, 11'b00000001000, 11'b00000000101, 11'b00000000000, 11'b11111111111, 11'b11111111101, 11'b11111111101, 11'b11111111101, 11'b11111111110, 11'b00000000010, 11'b11111111111, 11'b00000000000, 11'b00000000100, 11'b00000000000, 11'b00000000000, 11'b00000000000, 11'b00000001000, 11'b00000000001, 11'b00000000000, 11'b11111111100, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b00000000010}, 
{11'b11111111111, 11'b00000000000, 11'b11111111001, 11'b11111111101, 11'b00000001001, 11'b11111111111, 11'b11111111101, 11'b00000000111, 11'b11111111110, 11'b00000001001, 11'b00000000010, 11'b11111111100, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b11111111101, 11'b11111110111, 11'b00000001000, 11'b00000000100, 11'b00000010100, 11'b00000000110, 11'b00000000111, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b00000000001, 11'b00000000010, 11'b11111110010, 11'b11111111111, 11'b11111111111, 11'b11111111111}, 
{11'b00000000000, 11'b11111111101, 11'b11111111100, 11'b00000000000, 11'b11111111000, 11'b00000000000, 11'b00000000110, 11'b00000000011, 11'b00000000001, 11'b11111111100, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b11111111110, 11'b00000000110, 11'b11111111111, 11'b11111111111, 11'b11111110110, 11'b00000000000, 11'b11111111001, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b00000000000, 11'b00000000100, 11'b11111111101, 11'b11111111111, 11'b11111110001, 11'b00000000010}, 
{11'b00000001110, 11'b11111111111, 11'b00000000010, 11'b11111111100, 11'b11111111101, 11'b00000000001, 11'b00000000101, 11'b00000000000, 11'b00000010000, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b00000000011, 11'b11111111111, 11'b00000000001, 11'b00000000011, 11'b11111111111, 11'b11111110001, 11'b11111111110, 11'b11111111111, 11'b00000000011, 11'b00000000000, 11'b11111111111, 11'b00000000011, 11'b00000000000, 11'b11111110111, 11'b11111111100, 11'b00000000100, 11'b11111111111, 11'b00000001000, 11'b11111111111, 11'b11111111010}, 
{11'b00000000000, 11'b00000000011, 11'b11111111111, 11'b11111111110, 11'b11111110100, 11'b11111111111, 11'b00000000001, 11'b11111111110, 11'b00000000101, 11'b11111111110, 11'b11111111111, 11'b11111111110, 11'b11111111111, 11'b11111111110, 11'b00000000000, 11'b00000001010, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b00000000001, 11'b00000000100, 11'b00000000000, 11'b00000000000, 11'b00000000001, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b00000000000, 11'b00000000011}, 
{11'b11111110110, 11'b00000000100, 11'b00000000000, 11'b11111111100, 11'b11111110011, 11'b11111111111, 11'b00000000010, 11'b11111110011, 11'b00000010000, 11'b00000000010, 11'b00000000000, 11'b00000000011, 11'b00000000001, 11'b00000000000, 11'b00000001101, 11'b11111111101, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b11111110010, 11'b00000000000, 11'b00000000100, 11'b00000000001, 11'b00000000001, 11'b11111101010, 11'b11111110101, 11'b11111111000, 11'b00000000000, 11'b11111111111, 11'b00000001010, 11'b11111111001}, 
{11'b11111111111, 11'b11111111001, 11'b11111111100, 11'b11111110010, 11'b11111110111, 11'b00000001010, 11'b00000001001, 11'b11111111010, 11'b00000000001, 11'b11111111110, 11'b11111111100, 11'b11111110111, 11'b00000000011, 11'b11111110110, 11'b00000000110, 11'b11111111111, 11'b00000001010, 11'b11111111111, 11'b11111111111, 11'b11111111011, 11'b11111111110, 11'b11111111101, 11'b11111110111, 11'b00000000010, 11'b11111111111, 11'b11111111111, 11'b11111111000, 11'b00000001010, 11'b00000001000, 11'b11111111101, 11'b11111101011, 11'b00000000100}, 
{11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b11111111100, 11'b00000000000, 11'b00000000000, 11'b00000000010, 11'b00000000000, 11'b00000000011, 11'b11111111111, 11'b00000000000, 11'b00000000011, 11'b00000000000, 11'b00000000000, 11'b11111111011, 11'b11111111100, 11'b00000000000, 11'b00000000101, 11'b00000000001, 11'b00000000100, 11'b11111111111, 11'b11111111010, 11'b11111111111, 11'b00000000010, 11'b11111111111, 11'b00000000001, 11'b11111111111, 11'b00000000010, 11'b00000000000, 11'b00000000010, 11'b11111110011, 11'b11111111111}, 
{11'b00000001001, 11'b11111111111, 11'b00000000100, 11'b11111110110, 11'b11111111001, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b11111111011, 11'b00000000000, 11'b00000000000, 11'b00000000000, 11'b00000000000, 11'b11111111011, 11'b00000000100, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b00000000011, 11'b11111111001, 11'b00000000011, 11'b00000000100, 11'b00000000100, 11'b11111111111, 11'b00000010001, 11'b11111111011, 11'b00000001011, 11'b11111111110, 11'b11111110100, 11'b11111111010, 11'b00000000100}, 
{11'b11111101110, 11'b11111111111, 11'b11111111011, 11'b11111111111, 11'b00000001000, 11'b11111111010, 11'b11111111110, 11'b00000000111, 11'b00000000011, 11'b11111111000, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b00000000100, 11'b11111111000, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b11111111001, 11'b11111111111, 11'b00000000000, 11'b11111110101, 11'b00000000010, 11'b00000010011, 11'b00000001011, 11'b11111111110, 11'b11111111010, 11'b11111110001, 11'b00000000000, 11'b11111111110}, 
{11'b00000000000, 11'b00000000110, 11'b00000000000, 11'b11111111011, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b00000000110, 11'b00000000110, 11'b11111111011, 11'b00000000100, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b11111111010, 11'b00000001000, 11'b11111111110, 11'b11111110101, 11'b00000000011, 11'b11111111111, 11'b11111111111, 11'b00000000011, 11'b11111111101, 11'b11111111111, 11'b11111111110, 11'b00000000010, 11'b11111111011, 11'b00000000100, 11'b11111110100, 11'b00000000010, 11'b11111111111, 11'b00000000101}, 
{11'b11111111110, 11'b00000000000, 11'b00000000010, 11'b00000000000, 11'b11111111110, 11'b11111111111, 11'b00000000011, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b00000000000, 11'b00000000000, 11'b11111111100, 11'b00000000000, 11'b00000000011, 11'b00000000001, 11'b00000000011, 11'b11111111111, 11'b11111111111, 11'b00000000100, 11'b00000000111, 11'b11111111100, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b11111110001, 11'b11111111111, 11'b11111111101, 11'b11111111111, 11'b00000010010, 11'b00000000000, 11'b11111111001}, 
{11'b11111111111, 11'b11111111100, 11'b11111111111, 11'b00000000000, 11'b00000000010, 11'b11111111111, 11'b00000000000, 11'b11111111111, 11'b00000000010, 11'b11111111111, 11'b00000000000, 11'b00000000001, 11'b00000001001, 11'b11111111100, 11'b00000000000, 11'b11111100100, 11'b11111111111, 11'b11111111110, 11'b00000000000, 11'b11111111110, 11'b00000000010, 11'b11111111000, 11'b00000000011, 11'b00000000011, 11'b11111111111, 11'b11111101001, 11'b11111111000, 11'b11111111111, 11'b11111111111, 11'b00000001100, 11'b11111111111, 11'b00000000100}, 
{11'b00000000001, 11'b00000000000, 11'b00000000101, 11'b11111111100, 11'b11111111101, 11'b00000000111, 11'b11111111010, 11'b00000000001, 11'b11111110110, 11'b00000000000, 11'b00000000000, 11'b11111111101, 11'b00000000000, 11'b00000000000, 11'b11111111001, 11'b00000001101, 11'b11111111000, 11'b11111111111, 11'b00000000011, 11'b11111111111, 11'b00000000010, 11'b11111110000, 11'b00000001010, 11'b11111111111, 11'b11111111100, 11'b00000001111, 11'b00000000100, 11'b11111111010, 11'b11111111011, 11'b11111101110, 11'b11111111111, 11'b00000000000}, 
{11'b11111111111, 11'b00000000000, 11'b11111111110, 11'b11111110111, 11'b11111111111, 11'b11111110011, 11'b00000000000, 11'b00000001001, 11'b00000000111, 11'b00000000000, 11'b00000000000, 11'b11111111100, 11'b00000001010, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b00000001101, 11'b00000000000, 11'b11111111110, 11'b11111111110, 11'b11111110101, 11'b00000000100, 11'b00000000000, 11'b00000000000, 11'b00000000001, 11'b11111111101, 11'b11111110001, 11'b00000001000, 11'b11111110001, 11'b00000000001, 11'b11111111101, 11'b00000000000}, 
{11'b00000000001, 11'b00000000101, 11'b00000000000, 11'b11111111111, 11'b11111110001, 11'b00000000000, 11'b11111111111, 11'b00000000111, 11'b00000001000, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b00000000000, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b00000000101, 11'b11111111100, 11'b11111110010, 11'b11111111110, 11'b11111111100, 11'b11111111100, 11'b11111111101, 11'b11111111111, 11'b11111111101, 11'b11111111111, 11'b11111111111, 11'b00000000100, 11'b11111111111, 11'b00000001110}
};

localparam logic signed [10:0] bias [32] = '{
11'b00000101111,  // 1.474280834197998
11'b00000010110,  // 0.6914801001548767
11'b00000101110,  // 1.4406442642211914
11'b00000101101,  // 1.408045768737793
11'b00000011111,  // 0.9864811301231384
11'b00000011011,  // 0.8636202812194824
11'b11111101100,  // -0.6153604388237
11'b00000001111,  // 0.4839226007461548
11'b00000001111,  // 0.4862793982028961
11'b00000001011,  // 0.37162142992019653
11'b00000001110,  // 0.45989668369293213
11'b00000101001,  // 1.2998151779174805
11'b11111011111,  // -1.016528844833374
11'b11111110100,  // -0.35249894857406616
11'b00000001110,  // 0.44582197070121765
11'b11111111100,  // -0.1119980737566948
11'b11111111101,  // -0.06717441976070404
11'b00000000000,  // 0.00487547367811203
11'b00000000110,  // 0.1946917623281479
11'b11111100111,  // -0.7796769738197327
11'b00000010111,  // 0.7287401556968689
11'b00000110110,  // 1.714877724647522
11'b11111001100,  // -1.5971007347106934
11'b00000000010,  // 0.07393483817577362
11'b00000001010,  // 0.3225609362125397
11'b00000011011,  // 0.8453295230865479
11'b00000011100,  // 0.898597240447998
11'b00000001000,  // 0.2548799514770508
11'b00000011111,  // 0.9735668301582336
11'b00000100100,  // 1.1261906623840332
11'b00000001110,  // 0.44768181443214417
11'b11110110100   // -2.3676068782806396
};
endpackage