// Width: 15
// NFRAC: 7
package dense_1_15_7;

localparam logic signed [14:0] weights [16][64] = '{ 
{15'b000000000100000, 15'b111111110101100, 15'b111111111101000, 15'b111111111100011, 15'b111111111001100, 15'b000000000001110, 15'b111111101111011, 15'b000000000000000, 15'b000000000000111, 15'b000000000100001, 15'b000000000000000, 15'b111111111001100, 15'b111111111111111, 15'b000000000011010, 15'b000000000000100, 15'b111111111011110, 15'b000000000011101, 15'b000000000000111, 15'b000000000000000, 15'b111111111111111, 15'b000000000110000, 15'b111111111010101, 15'b111111111111101, 15'b000000000111100, 15'b111111111010110, 15'b111111110101000, 15'b111111111011100, 15'b111111111100111, 15'b111111111110010, 15'b111111111111111, 15'b000000000000100, 15'b000000000011111, 15'b000000000011001, 15'b111111111111110, 15'b000000000000000, 15'b000000000100111, 15'b111111111111101, 15'b111111111011111, 15'b000000000000011, 15'b000000000011000, 15'b111111111111110, 15'b000000000100011, 15'b111111111011101, 15'b000000001110110, 15'b111111111111111, 15'b000000000111001, 15'b000000000000000, 15'b000000000010111, 15'b000000000011001, 15'b111111111111100, 15'b000000000000000, 15'b000000000010100, 15'b000000000011011, 15'b000000000001001, 15'b111111111110001, 15'b111111111011000, 15'b000000001000100, 15'b111111111000000, 15'b000000000111011, 15'b111111111010010, 15'b000000001100101, 15'b111111111111111, 15'b000000000000001, 15'b000000000001010}, 
{15'b000000000000000, 15'b111111111010110, 15'b111111111101111, 15'b111111111011100, 15'b111111111010111, 15'b000000000001101, 15'b111111110011111, 15'b111111111111111, 15'b111111111100010, 15'b000000000010110, 15'b000000000000000, 15'b111111111110100, 15'b000000000011001, 15'b000000000000000, 15'b111111111111111, 15'b000000000011010, 15'b111111111111111, 15'b000000000000000, 15'b111111111101000, 15'b111111111011111, 15'b000000000111000, 15'b111111111110101, 15'b000000000000110, 15'b000000001011001, 15'b000000000100000, 15'b111111111100010, 15'b111111111100010, 15'b111111111111111, 15'b111111111110011, 15'b111111111001100, 15'b111111111111000, 15'b000000000111010, 15'b000000000100011, 15'b000000001000110, 15'b000000001010000, 15'b000000000000110, 15'b111111111110000, 15'b111111111001000, 15'b000000000000111, 15'b000000000011000, 15'b000000000000010, 15'b000000000011010, 15'b111111111100100, 15'b000000000100000, 15'b000000000010110, 15'b000000000000110, 15'b111111111010100, 15'b000000000001010, 15'b000000000100001, 15'b000000000000011, 15'b000000000000011, 15'b000000010010100, 15'b111111111110110, 15'b111111111110011, 15'b111111111111001, 15'b111111111111111, 15'b000000000100000, 15'b111111111010000, 15'b000000001111110, 15'b000000000000000, 15'b000000001000010, 15'b000000000011110, 15'b000000001101001, 15'b000000000010010}, 
{15'b111111111111111, 15'b000000000000000, 15'b111111111110101, 15'b111111111101001, 15'b111111111101000, 15'b000000000000101, 15'b000000010111101, 15'b111111111111111, 15'b111111101011101, 15'b111111111111111, 15'b111111111111111, 15'b111111111111101, 15'b111111111100010, 15'b000000000000000, 15'b111111111111110, 15'b000000000010101, 15'b000000001110011, 15'b111111111111111, 15'b000000000001001, 15'b000000000000000, 15'b000000000110100, 15'b111111110100011, 15'b000000001001001, 15'b111111110100100, 15'b000000001111001, 15'b111111111010011, 15'b111111111100000, 15'b111111110100100, 15'b000000010100011, 15'b000000000100011, 15'b000000000000001, 15'b000000001000010, 15'b000000010000010, 15'b111111101100111, 15'b111111111110011, 15'b000000000000100, 15'b111111111100010, 15'b000000001110010, 15'b111111111111010, 15'b000000000101000, 15'b000000000101010, 15'b000000000101111, 15'b111111111111111, 15'b111111111111111, 15'b111111111111101, 15'b000000000010100, 15'b111111111011100, 15'b111111111101010, 15'b111111111111101, 15'b000000000110010, 15'b111111111101001, 15'b000000000010011, 15'b111111111111111, 15'b000000000010001, 15'b111111111101001, 15'b111111111111111, 15'b111111111011000, 15'b111111110101010, 15'b111111111111111, 15'b000000000000000, 15'b000000011000101, 15'b000000000000001, 15'b111111111111111, 15'b111111111011000}, 
{15'b111111111000101, 15'b111111111010000, 15'b111111110100111, 15'b000000000100111, 15'b111111111010111, 15'b111111101010011, 15'b111111111110001, 15'b111111111011000, 15'b000000000011100, 15'b111111111111111, 15'b000000010100001, 15'b111111111110010, 15'b111111110011011, 15'b000000001001010, 15'b000000000000011, 15'b111111111111111, 15'b111111111000111, 15'b111111111111111, 15'b000000000000000, 15'b111111111100011, 15'b111111101101100, 15'b111111111110001, 15'b111111110100110, 15'b000000000011001, 15'b111111111001110, 15'b111111110001010, 15'b000000000101000, 15'b000000001011110, 15'b000000010100101, 15'b111111111000101, 15'b111111110110101, 15'b000000000001001, 15'b000000001000000, 15'b111111110010100, 15'b111111111010111, 15'b000000000000000, 15'b111111110100011, 15'b000000000011111, 15'b111111111000111, 15'b000000000001111, 15'b000000000111010, 15'b000000000010100, 15'b000000000000000, 15'b000000000000010, 15'b000000001000110, 15'b111111111100110, 15'b111111111111111, 15'b111111111010011, 15'b111111111111111, 15'b111111111110011, 15'b111111110110001, 15'b000000000001011, 15'b111111111111111, 15'b000000000011011, 15'b000000000101000, 15'b000000001010010, 15'b111111110000100, 15'b111111110001001, 15'b111111110100101, 15'b000000001101110, 15'b000000011011111, 15'b111111110001100, 15'b111111111111001, 15'b000000000110111}, 
{15'b000000000101011, 15'b111111110110000, 15'b111111111011110, 15'b111111111111111, 15'b111111111101100, 15'b000000000101011, 15'b000000000011000, 15'b111111111111111, 15'b111111110110011, 15'b111111111100001, 15'b111111111010000, 15'b000000000000110, 15'b000000000000000, 15'b000000000000000, 15'b111111111111010, 15'b000000000101101, 15'b000000000010001, 15'b111111111001101, 15'b000000000000011, 15'b000000000000001, 15'b000000000011010, 15'b111111111110000, 15'b000000000001001, 15'b111111111111101, 15'b000000010001000, 15'b111111111101000, 15'b111111111011100, 15'b111111111001100, 15'b000000000000000, 15'b000000000010101, 15'b000000000001110, 15'b000000000100011, 15'b111111111111110, 15'b000000000001001, 15'b000000000010000, 15'b111111111111111, 15'b000000000000000, 15'b000000001110000, 15'b111111111011011, 15'b111111111110110, 15'b000000000110111, 15'b000000000011111, 15'b111111111000001, 15'b000000000000000, 15'b111111101110111, 15'b111111111111111, 15'b111111111110000, 15'b000000000000001, 15'b111111111111111, 15'b111111111111100, 15'b111111111111111, 15'b000000000011000, 15'b111111111111111, 15'b000000000101000, 15'b111111111100111, 15'b111111110100001, 15'b111111111000100, 15'b111111110111110, 15'b111111110110001, 15'b000000001011111, 15'b000000010101111, 15'b000000001100101, 15'b000000000001111, 15'b111111111111111}, 
{15'b111111111000110, 15'b111111110101111, 15'b000000000000000, 15'b000000000100111, 15'b000000000100100, 15'b111111111100100, 15'b000000001001010, 15'b111111111111111, 15'b000000000011111, 15'b111111111111111, 15'b111111111111110, 15'b111111111110110, 15'b111111111101001, 15'b000000001001010, 15'b111111111110100, 15'b000000000000000, 15'b111111110110000, 15'b111111111010010, 15'b000000000000000, 15'b111111111111111, 15'b111111111111001, 15'b111111111010111, 15'b111111111010111, 15'b000000000111011, 15'b111111111010111, 15'b111111111111111, 15'b000000000100000, 15'b111111111110110, 15'b111111110001000, 15'b111111111111111, 15'b111111111110111, 15'b111111111111110, 15'b111111111111110, 15'b000000000000101, 15'b000000000010000, 15'b000000000101100, 15'b000000000000001, 15'b111111111110011, 15'b111111111011110, 15'b111111111111111, 15'b111111111101010, 15'b111111110111100, 15'b000000000110011, 15'b000000000000001, 15'b000000001001101, 15'b000000000000000, 15'b111111111111111, 15'b000000000001100, 15'b111111111001010, 15'b000000000011101, 15'b000000000000000, 15'b111111111110011, 15'b111111111010001, 15'b000000000110001, 15'b111111111111111, 15'b000000000101100, 15'b000000000011011, 15'b000000000011010, 15'b111111111111101, 15'b111111111111110, 15'b111111110011000, 15'b111111111101111, 15'b111111111111000, 15'b111111111111111}, 
{15'b111111111011011, 15'b111111111010101, 15'b111111111001000, 15'b111111111110111, 15'b111111111101110, 15'b000000000001101, 15'b111111110100110, 15'b111111111101100, 15'b111111111100011, 15'b111111111111111, 15'b111111111011011, 15'b000000000101100, 15'b000000000000100, 15'b000000000010001, 15'b000000000100111, 15'b000000000000000, 15'b000000001100110, 15'b000000000001011, 15'b000000000011111, 15'b000000000100010, 15'b111111111101011, 15'b000000000101110, 15'b111111111100000, 15'b111111110111111, 15'b000000000010110, 15'b000000001000010, 15'b111111111111111, 15'b000000000000110, 15'b111111110000110, 15'b000000000100100, 15'b000000000100010, 15'b111111111010000, 15'b000000000111100, 15'b000000001010101, 15'b000000000000000, 15'b000000000101011, 15'b111111111111111, 15'b000000000100100, 15'b000000000011001, 15'b000000000000000, 15'b111111111110000, 15'b111111111010001, 15'b000000000010010, 15'b000000000111101, 15'b000000001000010, 15'b111111111101010, 15'b111111111110101, 15'b111111111100111, 15'b111111111101110, 15'b000000000001111, 15'b000000000000000, 15'b000000000000100, 15'b000000000000000, 15'b000000000010111, 15'b111111111101001, 15'b000000001100010, 15'b000000000101101, 15'b111111111111100, 15'b000000000110001, 15'b000000000011011, 15'b111111100101111, 15'b111111110110110, 15'b111111111101001, 15'b111111111111110}, 
{15'b000000000000000, 15'b000000000011110, 15'b111111111111111, 15'b111111111111111, 15'b111111111010110, 15'b111111111111100, 15'b111111111011111, 15'b000000000000000, 15'b000000000000011, 15'b000000000110001, 15'b000000000000001, 15'b111111111001111, 15'b111111111110111, 15'b000000000000000, 15'b111111111111001, 15'b111111111000110, 15'b111111110010011, 15'b111111111111111, 15'b111111110110010, 15'b111111111000110, 15'b111111111001110, 15'b000000000101100, 15'b000000000000110, 15'b111111111101101, 15'b111111111001000, 15'b000000000010011, 15'b000000000000000, 15'b000000000111111, 15'b000000001100111, 15'b111111111111010, 15'b000000000000000, 15'b000000000011101, 15'b111111110101000, 15'b111111111010000, 15'b000000000000111, 15'b000000000001011, 15'b111111111011100, 15'b000000000011110, 15'b000000000010000, 15'b111111111101100, 15'b111111111001010, 15'b111111111111011, 15'b000000000000100, 15'b111111111101010, 15'b000000000000111, 15'b000000000011101, 15'b111111111110000, 15'b000000000000011, 15'b000000000000000, 15'b111111111100100, 15'b111111111001110, 15'b000000000110101, 15'b000000000010000, 15'b111111111101001, 15'b000000000010000, 15'b111111111111000, 15'b111111111000011, 15'b111111111101110, 15'b111111111111001, 15'b111111111110111, 15'b000000001101010, 15'b000000000011000, 15'b111111111111001, 15'b111111111111111}, 
{15'b000000000000001, 15'b000000001001011, 15'b111111110110101, 15'b111111111100010, 15'b000000000101001, 15'b111111111100101, 15'b000000010011011, 15'b111111111011011, 15'b111111111111111, 15'b000000000100101, 15'b000000000100000, 15'b111111111111111, 15'b111111111111001, 15'b111111111000010, 15'b000000000100100, 15'b000000000010100, 15'b111111111100111, 15'b111111111111111, 15'b000000000000000, 15'b000000000000000, 15'b000000000100001, 15'b111111111000101, 15'b000000000110010, 15'b000000001001110, 15'b111111111110100, 15'b111111111111111, 15'b111111111111101, 15'b111111111111111, 15'b000000001011110, 15'b000000000000000, 15'b111111111011101, 15'b000000000000000, 15'b000000000110001, 15'b111111110011000, 15'b111111110111010, 15'b000000000011001, 15'b000000000010001, 15'b111111110110110, 15'b111111111100111, 15'b111111111100100, 15'b000000000110011, 15'b000000000110010, 15'b000000000000000, 15'b111111111011101, 15'b000000000000000, 15'b000000000110010, 15'b111111111111000, 15'b111111111111111, 15'b000000000000001, 15'b000000000011111, 15'b111111111111000, 15'b111111111100111, 15'b000000000101100, 15'b111111111100100, 15'b000000000100011, 15'b000000001001010, 15'b000000000000101, 15'b000000000100001, 15'b111111111001100, 15'b111111111010001, 15'b000000001101010, 15'b111111111101111, 15'b000000000000101, 15'b111111111110100}, 
{15'b000000000000010, 15'b111111111000110, 15'b000000000101111, 15'b111111111011011, 15'b111111111111111, 15'b000000000011011, 15'b111111110110101, 15'b000000000011000, 15'b000000000111110, 15'b000000000010011, 15'b000000000101110, 15'b000000000101001, 15'b111111111011000, 15'b111111111110110, 15'b111111111111001, 15'b000000000000000, 15'b111111110000101, 15'b000000000101001, 15'b111111111111011, 15'b000000000000011, 15'b111111111010010, 15'b000000000001000, 15'b000000000010011, 15'b111111111111111, 15'b111111111000101, 15'b111111111111001, 15'b111111111110101, 15'b000000010011111, 15'b111111110101011, 15'b000000000001000, 15'b000000000001100, 15'b111111111111000, 15'b111111111100011, 15'b000000000001110, 15'b111111111110101, 15'b111111111101110, 15'b111111111101001, 15'b111111111100101, 15'b111111111111101, 15'b111111111011001, 15'b000000000101001, 15'b000000000001111, 15'b000000000111111, 15'b000000000001011, 15'b000000000000100, 15'b111111111011010, 15'b000000000000000, 15'b111111111111111, 15'b111111111111111, 15'b000000000011000, 15'b000000000010110, 15'b000000000100101, 15'b111111111111111, 15'b111111111011010, 15'b000000000000001, 15'b000000000000000, 15'b000000000101001, 15'b111111111100110, 15'b111111110111001, 15'b000000001000111, 15'b111111111011010, 15'b000000010010100, 15'b111111111111101, 15'b111111111010010}, 
{15'b111111110110110, 15'b111111111111111, 15'b111111111001011, 15'b000000000011101, 15'b000000000100001, 15'b111111111110010, 15'b000000001000010, 15'b111111111101010, 15'b111111111000010, 15'b111111111010001, 15'b111111111011111, 15'b111111111000011, 15'b111111111100010, 15'b000000000011001, 15'b000000000000000, 15'b000000000000000, 15'b000000001101011, 15'b111111111111010, 15'b111111111111111, 15'b000000000110100, 15'b000000000100101, 15'b111111110110101, 15'b111111111001111, 15'b000000000011000, 15'b111111111001000, 15'b111111111111101, 15'b111111111011110, 15'b111111111010101, 15'b111111111001000, 15'b000000000100110, 15'b000000000011101, 15'b111111111101100, 15'b111111111110110, 15'b111111110000011, 15'b111111111101001, 15'b000000000000110, 15'b111111111101111, 15'b111111111011010, 15'b111111111111111, 15'b000000000001111, 15'b111111111110000, 15'b111111111111111, 15'b111111111111011, 15'b111111110101010, 15'b000000000000000, 15'b000000000000000, 15'b000000000101011, 15'b111111111110000, 15'b000000000110110, 15'b111111111100111, 15'b000000000100100, 15'b111111111111111, 15'b000000000011100, 15'b111111111001101, 15'b111111111111111, 15'b000000001000001, 15'b000000000101000, 15'b000000000100101, 15'b000000000000011, 15'b111111111001100, 15'b111111111011001, 15'b111111110101000, 15'b111111111111111, 15'b000000000001101}, 
{15'b000000000100111, 15'b000000000000000, 15'b000000000010000, 15'b111111111111111, 15'b000000000010011, 15'b111111111101110, 15'b000000000011110, 15'b000000000000101, 15'b000000000010001, 15'b000000000101011, 15'b111111111011110, 15'b111111111111101, 15'b111111111111110, 15'b111111111111110, 15'b111111110101011, 15'b111111111011001, 15'b000000001010000, 15'b111111111111100, 15'b111111111111001, 15'b000000000000000, 15'b111111111001111, 15'b000000000000001, 15'b000000000100000, 15'b000000000000100, 15'b000000000000100, 15'b000000000101011, 15'b000000000000000, 15'b000000000000100, 15'b000000000000000, 15'b111111111111001, 15'b111111111100110, 15'b111111110101010, 15'b000000000100001, 15'b000000000101011, 15'b111111111111100, 15'b111111111100001, 15'b000000000000000, 15'b111111110101100, 15'b111111111111010, 15'b111111111111111, 15'b000000000011001, 15'b111111111101111, 15'b111111111111111, 15'b000000001101100, 15'b000000000111001, 15'b111111111111111, 15'b111111111111111, 15'b111111111111111, 15'b111111111100001, 15'b000000000010010, 15'b000000000010010, 15'b000000000010110, 15'b000000000010100, 15'b000000000110001, 15'b000000000101100, 15'b000000001010100, 15'b111111111101110, 15'b000000000110010, 15'b000000000010011, 15'b111111111010110, 15'b000000000001110, 15'b111111111001110, 15'b111111111000111, 15'b111111111000000}, 
{15'b000000000000000, 15'b000000000011101, 15'b111111111100111, 15'b000000000000000, 15'b111111111111001, 15'b111111111111011, 15'b111111110101011, 15'b111111111111111, 15'b000000000100000, 15'b000000000011111, 15'b000000000011110, 15'b111111111001101, 15'b111111111110100, 15'b000000000100100, 15'b111111111111111, 15'b000000000000000, 15'b111111110010100, 15'b111111111111111, 15'b000000000101111, 15'b000000000001001, 15'b000000000011110, 15'b111111111110001, 15'b000000000011111, 15'b000000000110011, 15'b111111111010010, 15'b111111111011100, 15'b111111111111111, 15'b111111111110101, 15'b000000000001000, 15'b000000000000000, 15'b111111111111111, 15'b000000000101000, 15'b111111110100000, 15'b000000000101110, 15'b000000001000000, 15'b000000000001110, 15'b000000000001110, 15'b111111111110010, 15'b000000000001110, 15'b111111111110010, 15'b111111111011111, 15'b111111111111001, 15'b000000000010101, 15'b000000001011001, 15'b111111110010011, 15'b111111111000110, 15'b000000000011000, 15'b111111111110011, 15'b000000000111001, 15'b111111111100001, 15'b111111111010101, 15'b111111111011100, 15'b111111111111111, 15'b000000000001111, 15'b111111111101011, 15'b111111110010100, 15'b111111111101101, 15'b111111111111110, 15'b000000000000101, 15'b111111110110001, 15'b000000010001111, 15'b111111110111010, 15'b000000001000101, 15'b000000000010011}, 
{15'b000000000001010, 15'b111111111100111, 15'b000000001010000, 15'b111111111011001, 15'b111111111000100, 15'b000000000001011, 15'b000000000100111, 15'b000000000100110, 15'b111111111101001, 15'b111111111101011, 15'b000000000000110, 15'b000000000011101, 15'b000000000011110, 15'b000000000000110, 15'b111111111100101, 15'b000000000010000, 15'b000000000111100, 15'b111111111111110, 15'b111111111011100, 15'b000000000000000, 15'b000000000001001, 15'b000000000000010, 15'b111111111011010, 15'b000000000001110, 15'b000000001100100, 15'b000000000000001, 15'b000000000010111, 15'b111111110011010, 15'b111111111110110, 15'b000000000000001, 15'b111111111100110, 15'b111111111011000, 15'b000000000111010, 15'b111111111111100, 15'b111111111111011, 15'b111111111011000, 15'b000000000010001, 15'b000000000100101, 15'b111111111111110, 15'b111111111111010, 15'b111111111101000, 15'b000000000011101, 15'b000000000000000, 15'b111111110101000, 15'b000000000100111, 15'b000000000110011, 15'b111111111111111, 15'b000000000000011, 15'b111111111001000, 15'b111111111110110, 15'b111111111111111, 15'b111111111010111, 15'b000000000000000, 15'b111111111101001, 15'b000000000000111, 15'b111111110010111, 15'b111111111111111, 15'b111111111111111, 15'b000000000100011, 15'b000000001001000, 15'b111111110100111, 15'b000000001000010, 15'b000000000000100, 15'b111111111110110}, 
{15'b000000000100100, 15'b000000010011110, 15'b000000000111111, 15'b000000000100100, 15'b111111111000010, 15'b111111111010111, 15'b111111010110011, 15'b111111111000101, 15'b000000000110011, 15'b111111111111111, 15'b000000000100101, 15'b000000001101110, 15'b000000000001000, 15'b000000000000000, 15'b111111111111101, 15'b000000000000000, 15'b111111111100111, 15'b111111111100110, 15'b000000000011101, 15'b111111110111111, 15'b111111110101010, 15'b111111111110010, 15'b111111110110101, 15'b000000000000011, 15'b111111011011100, 15'b000000001101000, 15'b000000001111110, 15'b000000001001101, 15'b111111100100000, 15'b111111111010111, 15'b111111110100111, 15'b111111110010100, 15'b111111010111100, 15'b000000001010110, 15'b111111111111010, 15'b000000000101000, 15'b000000000000011, 15'b111111101001000, 15'b000000000000000, 15'b000000000000000, 15'b000000000000100, 15'b000000010000010, 15'b111111111100101, 15'b111111110101101, 15'b000000001110010, 15'b111111111000111, 15'b111111111010110, 15'b111111111001101, 15'b000000000111101, 15'b000000001000100, 15'b111111111110111, 15'b111111111010011, 15'b111111111111111, 15'b111111111110001, 15'b000000000000000, 15'b111111111001111, 15'b000000001001101, 15'b000000010001010, 15'b000000001011011, 15'b111111110001011, 15'b111111000100110, 15'b000000001110001, 15'b000000000001011, 15'b000000000101000}, 
{15'b111111111100001, 15'b000000000101011, 15'b000000000101000, 15'b111111111111111, 15'b111111111010000, 15'b111111111110100, 15'b111111111001110, 15'b111111111111000, 15'b000000000010011, 15'b111111111110110, 15'b111111111111100, 15'b111111111111010, 15'b111111111111111, 15'b111111111101000, 15'b111111111111100, 15'b111111111110011, 15'b000000000101000, 15'b111111111111111, 15'b111111110101101, 15'b000000000111011, 15'b000000001001100, 15'b000000000110101, 15'b111111111010111, 15'b111111111101110, 15'b111111111010011, 15'b111111111011010, 15'b000000000011101, 15'b000000000011101, 15'b000000000011100, 15'b000000000101110, 15'b000000000000100, 15'b000000000110001, 15'b111111111111010, 15'b000000000000000, 15'b000000000100110, 15'b000000000010000, 15'b111111111110111, 15'b111111111111110, 15'b000000000000000, 15'b111111111011010, 15'b111111111100011, 15'b111111111110001, 15'b111111111010010, 15'b000000000111001, 15'b000000000000000, 15'b111111111111111, 15'b111111111110101, 15'b111111111101101, 15'b111111110011000, 15'b111111111111011, 15'b111111111100011, 15'b111111111101101, 15'b111111111110011, 15'b000000000100001, 15'b000000001010111, 15'b000000000010111, 15'b111111111111110, 15'b111111111010100, 15'b111111111111100, 15'b000000000000000, 15'b000000000101001, 15'b111111111111101, 15'b000000000000101, 15'b000000000000000}
};

localparam logic signed [14:0] bias [64] = '{
15'b111111111111011,  // -0.037350185215473175
15'b000000000100011,  // 0.27355897426605225
15'b111111111110000,  // -0.12378914654254913
15'b111111111110111,  // -0.064457006752491
15'b000000000000110,  // 0.05452875792980194
15'b000000000001110,  // 0.11671770364046097
15'b000000000010001,  // 0.13640816509723663
15'b000000000001001,  // 0.07482525706291199
15'b000000000000101,  // 0.04674031585454941
15'b111111111100110,  // -0.20146161317825317
15'b111111111110011,  // -0.09910125285387039
15'b000000000010011,  // 0.15104414522647858
15'b111111111110010,  // -0.10221704095602036
15'b111111111101101,  // -0.1461549550294876
15'b111111111110100,  // -0.08641516417264938
15'b000000000010101,  // 0.16613510251045227
15'b111111111110101,  // -0.0836295336484909
15'b111111111111000,  // -0.05756539851427078
15'b111111111111011,  // -0.03229188174009323
15'b111111111111100,  // -0.028388574719429016
15'b000000000010000,  // 0.1260243058204651
15'b111111111111011,  // -0.037064336240291595
15'b000000000011000,  // 0.19336333870887756
15'b000000000000010,  // 0.02124214917421341
15'b000000000111111,  // 0.4985624849796295
15'b000000000000010,  // 0.0158411655575037
15'b111111111110101,  // -0.08296407759189606
15'b000000000001110,  // 0.11056788265705109
15'b000000000000001,  // 0.01173810102045536
15'b111111111110010,  // -0.10843746364116669
15'b000000000100011,  // 0.27439257502555847
15'b000000000001011,  // 0.09199801832437515
15'b000000000100011,  // 0.27419957518577576
15'b000000000100010,  // 0.27063727378845215
15'b111111111100000,  // -0.24828937649726868
15'b000000000001010,  // 0.07818280160427094
15'b111111111111111,  // -0.005749030504375696
15'b000000000001101,  // 0.10850494354963303
15'b000000000010001,  // 0.13591453433036804
15'b111111111110000,  // -0.12088628858327866
15'b111111111111000,  // -0.05666546896100044
15'b000000000001011,  // 0.09311636537313461
15'b000000000000111,  // 0.05477767437696457
15'b000000000000011,  // 0.029585206881165504
15'b111111111011000,  // -0.31209176778793335
15'b111111111110101,  // -0.08465463668107986
15'b111111111101010,  // -0.16775836050510406
15'b000000000010010,  // 0.14762157201766968
15'b111111111100001,  // -0.23618532717227936
15'b000000000001000,  // 0.06535740196704865
15'b111111111101111,  // -0.12853026390075684
15'b111111111101110,  // -0.13802281022071838
15'b111111111101100,  // -0.15156887471675873
15'b000000000001010,  // 0.07979883998632431
15'b000000000010111,  // 0.18141601979732513
15'b111111111111001,  // -0.054039113223552704
15'b111111111111110,  // -0.010052933357656002
15'b000000000001000,  // 0.06611225008964539
15'b000000000000110,  // 0.05053366720676422
15'b000000000000011,  // 0.026860840618610382
15'b000000000000100,  // 0.03283466026186943
15'b000000000010011,  // 0.15558314323425293
15'b111111111011011,  // -0.2863388657569885
15'b111111111110100   // -0.08769102394580841
};
endpackage