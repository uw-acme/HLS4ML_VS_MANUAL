// Width: 13
// NFRAC: 6
package dense_3_13_6;

localparam logic signed [12:0] weights [32][32] = '{ 
{13'b1111111111100, 13'b1111111100100, 13'b1111111100110, 13'b1111111110011, 13'b0000000010101, 13'b0000000000010, 13'b1111111111111, 13'b1111111111111, 13'b1111111111111, 13'b1111111111111, 13'b0000000001000, 13'b1111111011110, 13'b1111111111100, 13'b0000000110110, 13'b1111111110000, 13'b1111111000100, 13'b1111111111101, 13'b0000000000111, 13'b0000000011011, 13'b1111111101001, 13'b1111110111011, 13'b1111111111101, 13'b0000000000011, 13'b1111111100110, 13'b0000000000000, 13'b0000001000000, 13'b1111110100010, 13'b1111111110001, 13'b1111111100111, 13'b1111111110110, 13'b0000000011011, 13'b1111111110101}, 
{13'b0000000101111, 13'b0000001101110, 13'b0000000011001, 13'b1111111010101, 13'b0000000001111, 13'b1111111101110, 13'b1111111111001, 13'b0000001000101, 13'b0000000000000, 13'b1111111111111, 13'b1111111111101, 13'b1111111011010, 13'b1111111110011, 13'b0000000100010, 13'b1111101111001, 13'b1111111100001, 13'b1111111111111, 13'b1111111111111, 13'b1111111111100, 13'b1111111110101, 13'b1111111101111, 13'b1111111101110, 13'b0000000000001, 13'b1111111111111, 13'b1111111111111, 13'b1111110111011, 13'b0000000000000, 13'b0000000011110, 13'b1111111111011, 13'b1111111010011, 13'b0000000000000, 13'b0000000000010}, 
{13'b1111111000000, 13'b0000000001011, 13'b0000000000000, 13'b0000000010100, 13'b1111111010111, 13'b0000000000000, 13'b0000000000000, 13'b1111111001010, 13'b0000000100010, 13'b1111111101111, 13'b1111111101111, 13'b1111110100000, 13'b1111111101100, 13'b0000000100000, 13'b0000000010000, 13'b1111111111111, 13'b1111111111000, 13'b1111111111110, 13'b1111111001011, 13'b0000000000000, 13'b0000000000111, 13'b0000000000100, 13'b0000000001101, 13'b0000000111000, 13'b0000000000010, 13'b1111111001101, 13'b0000000110001, 13'b0000000000000, 13'b0000000001010, 13'b1111111111110, 13'b0000000000000, 13'b0000010010001}, 
{13'b0000000110101, 13'b1111111111111, 13'b1111111110011, 13'b0000001010011, 13'b0000001001110, 13'b0000000000000, 13'b0000000000100, 13'b0000000110100, 13'b1111111100110, 13'b1111111111111, 13'b1111111001011, 13'b0000000000111, 13'b0000000010001, 13'b1111111010000, 13'b0000000000101, 13'b1111111110101, 13'b1111111111111, 13'b1111111101000, 13'b0000000000010, 13'b0000000000011, 13'b0000000000001, 13'b1111111111011, 13'b0000001001100, 13'b0000000101011, 13'b0000000101010, 13'b0000000011111, 13'b0000000101011, 13'b0000000000000, 13'b1111111111000, 13'b0000000111001, 13'b0000000011111, 13'b1111111110100}, 
{13'b0000001000000, 13'b1111111111010, 13'b1111111010011, 13'b1111110011111, 13'b0000000111101, 13'b0000000000000, 13'b1111111001011, 13'b1111111011011, 13'b1111111111010, 13'b1111110011000, 13'b1111101110010, 13'b0000000111100, 13'b0000001010101, 13'b0000001000010, 13'b1111110110110, 13'b1111110011100, 13'b0000000000000, 13'b1111111101101, 13'b0000000011001, 13'b0000000010001, 13'b1111111100111, 13'b1111111111111, 13'b0000001011100, 13'b1111101010000, 13'b0000000001011, 13'b1111110101011, 13'b0000000001000, 13'b1111111100000, 13'b1111111011001, 13'b1111111111111, 13'b0000000001000, 13'b0000001001010}, 
{13'b0000000000101, 13'b1111111111010, 13'b1111111011000, 13'b1111111011110, 13'b0000000101111, 13'b0000000000000, 13'b1111111011100, 13'b1111111101110, 13'b1111111001001, 13'b1111111110111, 13'b1111111111111, 13'b0000000010100, 13'b0000000000000, 13'b0000000101101, 13'b1111110111111, 13'b1111111101111, 13'b0000000001011, 13'b1111111011010, 13'b1111111100110, 13'b1111111111111, 13'b0000000000001, 13'b0000000100110, 13'b0000000111011, 13'b1111111111110, 13'b1111111111111, 13'b0000000110011, 13'b1111110111001, 13'b1111111111111, 13'b1111111100001, 13'b1111111111011, 13'b1111111111111, 13'b0000000000000}, 
{13'b0000000001000, 13'b1111111010101, 13'b0000000001101, 13'b1111111111011, 13'b1111111111111, 13'b0000000010011, 13'b1111111110010, 13'b1111110101001, 13'b1111111111111, 13'b1111111100101, 13'b1111111000101, 13'b0000000111100, 13'b0000000000000, 13'b0000001010111, 13'b0000001101010, 13'b0000000000000, 13'b1111111111111, 13'b1111111010111, 13'b1111111111000, 13'b0000000100010, 13'b1111110011111, 13'b0000000010011, 13'b0000000101001, 13'b0000000000010, 13'b0000000010011, 13'b0000010011111, 13'b1111111001101, 13'b1111111110100, 13'b1111111100111, 13'b0000000111110, 13'b1111111111001, 13'b1111111101010}, 
{13'b1111110110011, 13'b0000000000011, 13'b1111110101111, 13'b0000000110111, 13'b0000010000011, 13'b0000000001110, 13'b0000000000000, 13'b0000000000110, 13'b1111111111111, 13'b0000000010000, 13'b0000010100110, 13'b1111111111111, 13'b0000000110000, 13'b0000001001111, 13'b0000001100010, 13'b0000010000110, 13'b0000000000000, 13'b1111111000010, 13'b0000000101011, 13'b1111111111111, 13'b1111110101110, 13'b1111111100010, 13'b0000000000001, 13'b1111111110101, 13'b1111110111111, 13'b0000011110000, 13'b1111111100011, 13'b0000000000000, 13'b0000000000000, 13'b0000001110001, 13'b0000000001011, 13'b0000000110010}, 
{13'b0000000110110, 13'b1111111111101, 13'b0000000000000, 13'b1111111111010, 13'b0000000001010, 13'b1111111111011, 13'b1111111111111, 13'b0000000010100, 13'b0000000011011, 13'b1111111011100, 13'b0000000010001, 13'b0000000010111, 13'b0000000000001, 13'b0000000101010, 13'b1111111100011, 13'b1111110011001, 13'b0000000000000, 13'b1111111111110, 13'b1111111111100, 13'b1111111000000, 13'b1111111111111, 13'b0000000000000, 13'b1111111100110, 13'b1111111111110, 13'b1111111110011, 13'b0000000010011, 13'b0000000101111, 13'b1111111110000, 13'b1111111111001, 13'b1111111111010, 13'b0000000000011, 13'b1111111001101}, 
{13'b1111111101001, 13'b0000000110001, 13'b0000000000000, 13'b0000000000000, 13'b0000001100101, 13'b0000000101001, 13'b1111111111111, 13'b1111110111000, 13'b0000000001111, 13'b1111110100110, 13'b1111101001100, 13'b1111111111111, 13'b0000000000000, 13'b0000000110110, 13'b0000000001110, 13'b0000000000000, 13'b1111111010101, 13'b0000000000000, 13'b0000000000000, 13'b0000000000111, 13'b0000000011111, 13'b1111111111100, 13'b1111111010001, 13'b0000000000001, 13'b1111111111110, 13'b0000010001010, 13'b0000000101001, 13'b1111111111111, 13'b1111111110110, 13'b0000001010101, 13'b1111111111010, 13'b1111111110100}, 
{13'b1111110111101, 13'b0000000010110, 13'b1111111111011, 13'b1111111111111, 13'b1111111100000, 13'b1111111001111, 13'b0000000000110, 13'b0000000010010, 13'b1111111111111, 13'b1111111101010, 13'b1111110110110, 13'b0000000011001, 13'b0000000100110, 13'b0000000000000, 13'b0000001101011, 13'b1111110111000, 13'b0000000001101, 13'b1111111001101, 13'b0000000100100, 13'b1111111111111, 13'b1111111111011, 13'b0000000001000, 13'b0000000001111, 13'b0000000000000, 13'b1111111000000, 13'b0000000000011, 13'b1111110111000, 13'b1111111111010, 13'b1111111111111, 13'b0000001010110, 13'b1111111100111, 13'b0000000000000}, 
{13'b1111111111111, 13'b0000000001110, 13'b0000000000000, 13'b0000000110010, 13'b1111111110001, 13'b1111111111010, 13'b0000000000111, 13'b1111111111111, 13'b1111111111010, 13'b0000001010010, 13'b0000001011001, 13'b0000000000000, 13'b1111111010101, 13'b1111110100110, 13'b1111111111001, 13'b0000000000000, 13'b0000000000000, 13'b1111111110111, 13'b1111111000011, 13'b0000000110000, 13'b0000000000000, 13'b0000000101111, 13'b1111111111111, 13'b0000001000111, 13'b0000000001111, 13'b0000000100111, 13'b0000000111010, 13'b1111111111001, 13'b1111111001101, 13'b1111111000111, 13'b1111111111111, 13'b1111110101010}, 
{13'b1111111100011, 13'b1111111111111, 13'b0000000001111, 13'b1111111001010, 13'b0000000001011, 13'b1111111111111, 13'b1111111100100, 13'b1111111111110, 13'b1111111101111, 13'b0000000000100, 13'b0000000001001, 13'b1111111110110, 13'b0000000000010, 13'b0000000011000, 13'b1111110101111, 13'b1111111100000, 13'b0000000011101, 13'b1111111101001, 13'b0000000000000, 13'b1111111111100, 13'b0000000011000, 13'b0000000000001, 13'b1111111111100, 13'b0000000000101, 13'b0000000100010, 13'b1111111110010, 13'b0000000000000, 13'b1111111000110, 13'b1111111100110, 13'b1111111111111, 13'b0000000010110, 13'b0000000000000}, 
{13'b1111110111101, 13'b0000000110101, 13'b1111111111111, 13'b1111111111111, 13'b1111111111110, 13'b0000000010110, 13'b1111111111111, 13'b0000001100010, 13'b1111111111110, 13'b1111111111111, 13'b0000000011010, 13'b0000000000101, 13'b0000000000000, 13'b0000000000000, 13'b0000000001111, 13'b0000000101010, 13'b0000000010110, 13'b0000000010101, 13'b1111111111110, 13'b0000000100111, 13'b0000000001100, 13'b0000000000101, 13'b1111111111110, 13'b0000000100000, 13'b1111111110011, 13'b1111111010100, 13'b1111111110100, 13'b1111111111111, 13'b0000000001101, 13'b0000000000011, 13'b0000000011001, 13'b0000000111101}, 
{13'b1111111111101, 13'b1111111001110, 13'b0000000000110, 13'b1111111111111, 13'b0000001110101, 13'b1111111100101, 13'b1111110110110, 13'b0000000000000, 13'b0000000000000, 13'b1111111111100, 13'b0000000000110, 13'b0000000110111, 13'b0000000101001, 13'b0000000000001, 13'b0000000000100, 13'b1111111101001, 13'b0000000000100, 13'b1111111111011, 13'b0000000000000, 13'b0000000001001, 13'b1111111111011, 13'b0000000000010, 13'b0000000100010, 13'b0000000000100, 13'b1111111111110, 13'b1111111001011, 13'b0000000011010, 13'b1111111111111, 13'b1111111111111, 13'b1111111110010, 13'b1111111111101, 13'b1111111110111}, 
{13'b0000000000000, 13'b1111111110111, 13'b1111111101111, 13'b1111111100100, 13'b1111110111010, 13'b0000001001110, 13'b0000000000000, 13'b0000000010101, 13'b0000000100100, 13'b0000000000001, 13'b1111111111011, 13'b0000000111100, 13'b0000000011100, 13'b1111111010001, 13'b1111111101011, 13'b1111111111010, 13'b1111111001101, 13'b1111111111101, 13'b0000000000000, 13'b1111111111111, 13'b0000000010011, 13'b1111111101110, 13'b0000000000000, 13'b0000000001001, 13'b1111111111111, 13'b1111111010100, 13'b0000000010100, 13'b0000000000000, 13'b0000000000101, 13'b0000000000001, 13'b1111111010111, 13'b0000000000010}, 
{13'b1111111100110, 13'b1111111101011, 13'b0000000001001, 13'b1111111110000, 13'b1111111110100, 13'b0000000001110, 13'b1111111111111, 13'b0000000000100, 13'b0000000010000, 13'b1111111111111, 13'b0000000001111, 13'b1111111101111, 13'b1111111111110, 13'b1111111111111, 13'b0000000001101, 13'b1111111111111, 13'b0000000111110, 13'b1111111111101, 13'b0000000011111, 13'b1111111101010, 13'b0000000010100, 13'b0000000001000, 13'b0000000001010, 13'b0000000000100, 13'b1111111110101, 13'b1111111011100, 13'b1111111011110, 13'b0000000001101, 13'b1111111110101, 13'b0000000000000, 13'b1111111111100, 13'b0000000011101}, 
{13'b1111111111111, 13'b1111111001100, 13'b1111111001101, 13'b1111111111111, 13'b0000001010000, 13'b1111111110100, 13'b0000000000000, 13'b0000000111101, 13'b1111111101101, 13'b0000000000000, 13'b1111111001010, 13'b1111111000001, 13'b0000000111001, 13'b0000000010011, 13'b1111111110000, 13'b1111111011100, 13'b0000000010110, 13'b0000000000000, 13'b1111111100001, 13'b0000000000011, 13'b0000000001000, 13'b1111111110100, 13'b0000000100100, 13'b1111110000010, 13'b0000000000101, 13'b0000000011110, 13'b1111111111010, 13'b0000000000001, 13'b1111111100010, 13'b1111111111111, 13'b1111111100110, 13'b1111111111100}, 
{13'b0000000011011, 13'b0000000101100, 13'b0000001000110, 13'b1111111100101, 13'b0000000110101, 13'b0000000100111, 13'b0000000000000, 13'b0000000111010, 13'b0000000101101, 13'b1111111110010, 13'b0000001011001, 13'b1111111010011, 13'b0000001001111, 13'b0000000111001, 13'b1111101110110, 13'b1111111111111, 13'b0000000000000, 13'b0000000000000, 13'b0000000100001, 13'b1111110111111, 13'b0000000011100, 13'b1111111100100, 13'b1111111000001, 13'b1111111101011, 13'b0000000101010, 13'b1111110101011, 13'b1111111010101, 13'b1111111111010, 13'b1111111111111, 13'b1111110110111, 13'b0000000110010, 13'b0000000000000}, 
{13'b1111111111001, 13'b0000000000000, 13'b1111111111111, 13'b1111111111111, 13'b1111111010011, 13'b0000000000001, 13'b0000000000001, 13'b1111111111110, 13'b1111111111100, 13'b1111111111010, 13'b0000000010001, 13'b1111111111111, 13'b0000000001010, 13'b1111111010100, 13'b0000000001101, 13'b1111111111111, 13'b0000000010010, 13'b0000000111001, 13'b1111111010010, 13'b0000000000110, 13'b1111111110011, 13'b0000000010000, 13'b0000000011000, 13'b1111111110101, 13'b1111111011111, 13'b0000000000010, 13'b0000001101010, 13'b1111111111100, 13'b1111111111110, 13'b0000000101001, 13'b0000000000000, 13'b0000001101110}, 
{13'b1111110111101, 13'b0000000000100, 13'b1111111100100, 13'b0000000110001, 13'b0000000001110, 13'b1111111111011, 13'b1111111111111, 13'b1111111111111, 13'b1111111011001, 13'b1111111111011, 13'b0000000000000, 13'b1111110111000, 13'b0000000000001, 13'b1111111111010, 13'b1111111111111, 13'b1111111111111, 13'b1111111110001, 13'b0000000000000, 13'b0000000000000, 13'b0000000010100, 13'b0000000000010, 13'b0000000000000, 13'b0000000000000, 13'b1111111111110, 13'b0000000000000, 13'b0000000000010, 13'b0000001001010, 13'b1111111111111, 13'b1111111111111, 13'b1111111111010, 13'b0000000010110, 13'b1111111111100}, 
{13'b1111111111111, 13'b1111111101100, 13'b0000000011010, 13'b0000000000101, 13'b1111111010000, 13'b0000000000000, 13'b0000000100100, 13'b1111111111111, 13'b0000000000000, 13'b1111111110011, 13'b0000000001110, 13'b0000000000010, 13'b0000000101001, 13'b1111110111001, 13'b1111111110011, 13'b1111111111101, 13'b0000000011011, 13'b1111111001110, 13'b0000000000010, 13'b1111110011111, 13'b1111111111101, 13'b1111111110000, 13'b1111111111010, 13'b0000000100101, 13'b1111111110110, 13'b1111111011100, 13'b0000000001011, 13'b0000000000000, 13'b0000000110010, 13'b0000001000010, 13'b1111111010110, 13'b1111111000110}, 
{13'b0000000001000, 13'b0000000000011, 13'b1111111001010, 13'b1111111111000, 13'b1111111111111, 13'b0000000000000, 13'b0000000001101, 13'b0000000110100, 13'b0000000000000, 13'b0000000000010, 13'b0000000001000, 13'b1111110111010, 13'b1111111110111, 13'b1111110110010, 13'b0000000111101, 13'b0000000000000, 13'b1111111111111, 13'b1111110101101, 13'b1111111111111, 13'b1111111110110, 13'b1111111111101, 13'b0000000000000, 13'b0000000000111, 13'b1111111101100, 13'b0000000000110, 13'b0000000110100, 13'b0000000110110, 13'b0000000110001, 13'b0000000100111, 13'b0000000000000, 13'b0000000001110, 13'b0000001100100}, 
{13'b1111111111100, 13'b1111111100001, 13'b0000000110001, 13'b1111111110010, 13'b0000000001000, 13'b0000000010101, 13'b1111111111111, 13'b1111111011011, 13'b1111111110101, 13'b1111110110011, 13'b0000000111001, 13'b0000000000000, 13'b0000000110101, 13'b0000001010101, 13'b1111111110001, 13'b1111110010000, 13'b1111111110010, 13'b0000000111100, 13'b1111111011011, 13'b1111111100101, 13'b0000000000111, 13'b0000000000000, 13'b1111110111010, 13'b1111111100111, 13'b1111111111010, 13'b1111111110000, 13'b0000000001110, 13'b0000001011010, 13'b0000000011111, 13'b1111111111111, 13'b0000000001010, 13'b0000000000011}, 
{13'b0000000000101, 13'b0000000111010, 13'b0000000000000, 13'b0000000100101, 13'b0000001101010, 13'b1111111101010, 13'b1111111111111, 13'b1111111111010, 13'b0000000100101, 13'b1111111100111, 13'b1111111111111, 13'b0000000101010, 13'b0000000000001, 13'b0000000000011, 13'b1111100111100, 13'b1111111110101, 13'b0000000000000, 13'b0000000011001, 13'b1111111111111, 13'b0000000100110, 13'b1111111111111, 13'b1111111101001, 13'b1111110111000, 13'b0000000010000, 13'b0000000100100, 13'b1111101110010, 13'b1111111111111, 13'b0000000000000, 13'b0000001000101, 13'b1111110011001, 13'b0000000000000, 13'b1111111111111}, 
{13'b0000000000001, 13'b1111111010100, 13'b0000000000110, 13'b1111111111110, 13'b0000000000110, 13'b0000001000011, 13'b1111110100011, 13'b0000000000100, 13'b0000000110110, 13'b1111111010100, 13'b1111111111101, 13'b0000000000110, 13'b1111111111110, 13'b0000000010110, 13'b0000000001101, 13'b1111111111101, 13'b0000000001000, 13'b0000000000000, 13'b0000000000010, 13'b0000000110000, 13'b1111111111100, 13'b1111111000010, 13'b1111110110010, 13'b1111111100111, 13'b1111110110100, 13'b0000000011010, 13'b0000001001111, 13'b0000000101111, 13'b1111111111110, 13'b1111111010000, 13'b1111111011000, 13'b0000000000111}, 
{13'b0000000000110, 13'b1111111000010, 13'b1111111111101, 13'b0000000010011, 13'b1111111000010, 13'b0000000010101, 13'b1111111111111, 13'b1111111111111, 13'b1111111111111, 13'b0000000000000, 13'b0000000100001, 13'b1111111111101, 13'b0000000000001, 13'b0000000000000, 13'b0000000010000, 13'b1111111111101, 13'b0000000000000, 13'b1111111111111, 13'b1111111010110, 13'b1111110111111, 13'b1111111111111, 13'b1111110111011, 13'b1111111011001, 13'b1111111010000, 13'b0000001110001, 13'b0000000000010, 13'b1111111111010, 13'b0000000101000, 13'b0000001110010, 13'b0000000110010, 13'b1111101111000, 13'b1111111101000}, 
{13'b0000000110000, 13'b1111111111111, 13'b0000000100000, 13'b1111111111101, 13'b0000000111101, 13'b1111111101101, 13'b0000000001001, 13'b0000000110101, 13'b0000000100010, 13'b1111110111101, 13'b1111111111000, 13'b0000000001111, 13'b0000000001000, 13'b1111111111110, 13'b0000000001010, 13'b0000000000000, 13'b0000000101110, 13'b0000000000100, 13'b0000000101111, 13'b1111111110111, 13'b1111111101111, 13'b1111111110110, 13'b1111111111111, 13'b0000000100110, 13'b1111111100110, 13'b1111111111111, 13'b0000000000000, 13'b0000000000000, 13'b0000000000000, 13'b0000000100101, 13'b1111111010110, 13'b1111111111101}, 
{13'b1111111111111, 13'b1111111111100, 13'b1111111000100, 13'b0000000100100, 13'b0000000011100, 13'b1111111110001, 13'b1111111111111, 13'b1111111100010, 13'b0000000000000, 13'b1111111111111, 13'b1111111011001, 13'b1111111100000, 13'b0000000111101, 13'b0000000000000, 13'b1111111101111, 13'b1111111111111, 13'b0000000011011, 13'b1111111111111, 13'b1111111111111, 13'b1111111100100, 13'b0000000101000, 13'b0000000000000, 13'b0000000010011, 13'b1111111111100, 13'b0000000010100, 13'b0000000000000, 13'b0000000000000, 13'b0000000011110, 13'b1111111100111, 13'b1111111111010, 13'b0000000010100, 13'b1111111110010}, 
{13'b1111111111101, 13'b1111111011000, 13'b0000001001100, 13'b1111111110111, 13'b0000000011001, 13'b1111111011011, 13'b0000000000000, 13'b0000000000100, 13'b1111111000010, 13'b1111111111110, 13'b1111111110000, 13'b0000000000111, 13'b1111111010110, 13'b0000000010001, 13'b0000000011001, 13'b0000000001110, 13'b0000000001010, 13'b1111111111011, 13'b1111110100101, 13'b1111111111110, 13'b1111111111000, 13'b0000000010001, 13'b1111111110001, 13'b1111111111111, 13'b0000000011001, 13'b1111111111010, 13'b1111111111110, 13'b0000000110001, 13'b1111111001101, 13'b1111111011010, 13'b0000000101100, 13'b0000000000100}, 
{13'b0000000110111, 13'b0000000011001, 13'b0000000000000, 13'b1111111101011, 13'b1111111110101, 13'b1111111111111, 13'b0000000000000, 13'b1111111110111, 13'b1111111110000, 13'b1111111110000, 13'b0000000000000, 13'b0000000010100, 13'b0000000000000, 13'b0000000000110, 13'b1111111111010, 13'b0000000000000, 13'b1111111101100, 13'b0000000000000, 13'b1111111111101, 13'b1111111111111, 13'b0000000000000, 13'b0000000000111, 13'b0000000001100, 13'b0000000000000, 13'b0000000000000, 13'b1111110110001, 13'b1111111100110, 13'b0000000000000, 13'b0000000000010, 13'b0000000000000, 13'b1111111101001, 13'b0000000000010}, 
{13'b0000000011000, 13'b1111101111010, 13'b1111111111111, 13'b1111111110110, 13'b1111111100010, 13'b1111111111110, 13'b0000000000000, 13'b0000001000110, 13'b1111111111010, 13'b1111111111101, 13'b0000000001010, 13'b1111110101011, 13'b0000000000011, 13'b1111111000111, 13'b0000001011100, 13'b1111111111001, 13'b1111111100011, 13'b1111110111001, 13'b1111111111110, 13'b1111110100101, 13'b1111110011000, 13'b1111111111111, 13'b0000000000000, 13'b0000000000000, 13'b0000000011111, 13'b1111111111110, 13'b1111111011001, 13'b1111111110110, 13'b1111111111101, 13'b0000000000000, 13'b1111111111011, 13'b1111110100110}
};

localparam logic signed [12:0] bias [32] = '{
13'b0000000100001,  // 0.5280959606170654
13'b0000000110101,  // 0.8414360880851746
13'b0000000011001,  // 0.397830605506897
13'b0000000011010,  // 0.4105983078479767
13'b1111100010101,  // -3.657735586166382
13'b1111111000110,  // -0.8977976441383362
13'b0000001101101,  // 1.7051936388015747
13'b1111110101110,  // -1.2765135765075684
13'b1111111011010,  // -0.5837795734405518
13'b0000010101100,  // 2.699671983718872
13'b0000000001101,  // 0.2170683741569519
13'b0000000111000,  // 0.8814588785171509
13'b1111101010111,  // -2.634300947189331
13'b1111110000111,  // -1.877297282218933
13'b0000001101010,  // 1.6625694036483765
13'b0000010101111,  // 2.7459704875946045
13'b1111111100001,  // -0.47838035225868225
13'b0000001101100,  // 1.6984987258911133
13'b0000000110110,  // 0.8548859357833862
13'b0000001000000,  // 1.0045719146728516
13'b0000001011010,  // 1.4197649955749512
13'b0000000110101,  // 0.832463800907135
13'b0000000100010,  // 0.5434179306030273
13'b0000000111011,  // 0.9277304410934448
13'b1111111101010,  // -0.3426123857498169
13'b1111111011100,  // -0.5587119460105896
13'b1111111011000,  // -0.6208624839782715
13'b1111110101110,  // -1.2802538871765137
13'b0000000000011,  // 0.05940237268805504
13'b1111111001011,  // -0.8213341236114502
13'b0000000111000,  // 0.8783953189849854
13'b1111111000011   // -0.949700653553009
};
endpackage