// Width: 16
// NFRAC: 8
package dense_3_16_8;

localparam logic signed [15:0] weights [32][32] = '{ 
{16'b1111111111110011, 16'b1111111110010000, 16'b1111111110011000, 16'b1111111111001111, 16'b0000000001010111, 16'b0000000000001011, 16'b1111111111111100, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000100000, 16'b1111111101111001, 16'b1111111111110000, 16'b0000000011011000, 16'b1111111111000010, 16'b1111111100010001, 16'b1111111111110110, 16'b0000000000011100, 16'b0000000001101111, 16'b1111111110100110, 16'b1111111011101111, 16'b1111111111110100, 16'b0000000000001100, 16'b1111111110011000, 16'b0000000000000000, 16'b0000000100000011, 16'b1111111010001011, 16'b1111111111000111, 16'b1111111110011100, 16'b1111111111011001, 16'b0000000001101100, 16'b1111111111010111}, 
{16'b0000000010111111, 16'b0000000110111010, 16'b0000000001100110, 16'b1111111101010111, 16'b0000000000111110, 16'b1111111110111010, 16'b1111111111100100, 16'b0000000100010111, 16'b0000000000000001, 16'b1111111111111111, 16'b1111111111110111, 16'b1111111101101001, 16'b1111111111001100, 16'b0000000010001010, 16'b1111110111100100, 16'b1111111110000111, 16'b1111111111111111, 16'b1111111111111101, 16'b1111111111110010, 16'b1111111111010101, 16'b1111111110111101, 16'b1111111110111001, 16'b0000000000000100, 16'b1111111111111111, 16'b1111111111111110, 16'b1111111011101101, 16'b0000000000000011, 16'b0000000001111000, 16'b1111111111101111, 16'b1111111101001111, 16'b0000000000000000, 16'b0000000000001001}, 
{16'b1111111100000011, 16'b0000000000101111, 16'b0000000000000010, 16'b0000000001010010, 16'b1111111101011110, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111100101001, 16'b0000000010001001, 16'b1111111110111100, 16'b1111111110111101, 16'b1111111010000011, 16'b1111111110110000, 16'b0000000010000010, 16'b0000000001000011, 16'b1111111111111111, 16'b1111111111100010, 16'b1111111111111001, 16'b1111111100101111, 16'b0000000000000000, 16'b0000000000011111, 16'b0000000000010001, 16'b0000000000110101, 16'b0000000011100001, 16'b0000000000001001, 16'b1111111100110110, 16'b0000000011000100, 16'b0000000000000000, 16'b0000000000101010, 16'b1111111111111010, 16'b0000000000000000, 16'b0000001001000100}, 
{16'b0000000011010110, 16'b1111111111111111, 16'b1111111111001110, 16'b0000000101001111, 16'b0000000100111010, 16'b0000000000000000, 16'b0000000000010010, 16'b0000000011010000, 16'b1111111110011010, 16'b1111111111111111, 16'b1111111100101101, 16'b0000000000011110, 16'b0000000001000100, 16'b1111111101000000, 16'b0000000000010111, 16'b1111111111010111, 16'b1111111111111111, 16'b1111111110100010, 16'b0000000000001001, 16'b0000000000001110, 16'b0000000000000100, 16'b1111111111101101, 16'b0000000100110001, 16'b0000000010101111, 16'b0000000010101000, 16'b0000000001111111, 16'b0000000010101110, 16'b0000000000000000, 16'b1111111111100001, 16'b0000000011100111, 16'b0000000001111111, 16'b1111111111010011}, 
{16'b0000000100000000, 16'b1111111111101000, 16'b1111111101001110, 16'b1111111001111111, 16'b0000000011110100, 16'b0000000000000000, 16'b1111111100101101, 16'b1111111101101111, 16'b1111111111101000, 16'b1111111001100001, 16'b1111110111001010, 16'b0000000011110010, 16'b0000000101010110, 16'b0000000100001011, 16'b1111111011011001, 16'b1111111001110011, 16'b0000000000000000, 16'b1111111110110111, 16'b0000000001100110, 16'b0000000001000111, 16'b1111111110011111, 16'b1111111111111100, 16'b0000000101110001, 16'b1111110101000000, 16'b0000000000101101, 16'b1111111010101110, 16'b0000000000100001, 16'b1111111110000000, 16'b1111111101100111, 16'b1111111111111111, 16'b0000000000100011, 16'b0000000100101001}, 
{16'b0000000000010110, 16'b1111111111101010, 16'b1111111101100010, 16'b1111111101111010, 16'b0000000010111110, 16'b0000000000000000, 16'b1111111101110000, 16'b1111111110111010, 16'b1111111100100100, 16'b1111111111011111, 16'b1111111111111111, 16'b0000000001010010, 16'b0000000000000000, 16'b0000000010110111, 16'b1111111011111101, 16'b1111111110111110, 16'b0000000000101101, 16'b1111111101101001, 16'b1111111110011010, 16'b1111111111111111, 16'b0000000000000110, 16'b0000000010011001, 16'b0000000011101111, 16'b1111111111111010, 16'b1111111111111111, 16'b0000000011001101, 16'b1111111011100110, 16'b1111111111111111, 16'b1111111110000110, 16'b1111111111101101, 16'b1111111111111110, 16'b0000000000000011}, 
{16'b0000000000100001, 16'b1111111101010101, 16'b0000000000110111, 16'b1111111111101100, 16'b1111111111111100, 16'b0000000001001101, 16'b1111111111001001, 16'b1111111010100101, 16'b1111111111111111, 16'b1111111110010101, 16'b1111111100010110, 16'b0000000011110001, 16'b0000000000000011, 16'b0000000101011110, 16'b0000000110101000, 16'b0000000000000001, 16'b1111111111111111, 16'b1111111101011110, 16'b1111111111100000, 16'b0000000010001011, 16'b1111111001111111, 16'b0000000001001111, 16'b0000000010100111, 16'b0000000000001001, 16'b0000000001001100, 16'b0000001001111100, 16'b1111111100110110, 16'b1111111111010001, 16'b1111111110011110, 16'b0000000011111001, 16'b1111111111100110, 16'b1111111110101001}, 
{16'b1111111011001110, 16'b0000000000001100, 16'b1111111010111101, 16'b0000000011011110, 16'b0000001000001110, 16'b0000000000111011, 16'b0000000000000001, 16'b0000000000011000, 16'b1111111111111111, 16'b0000000001000001, 16'b0000001010011010, 16'b1111111111111111, 16'b0000000011000011, 16'b0000000100111110, 16'b0000000110001001, 16'b0000001000011001, 16'b0000000000000000, 16'b1111111100001011, 16'b0000000010101100, 16'b1111111111111101, 16'b1111111010111001, 16'b1111111110001011, 16'b0000000000000110, 16'b1111111111010101, 16'b1111111011111111, 16'b0000001111000000, 16'b1111111110001111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000111000100, 16'b0000000000101101, 16'b0000000011001000}, 
{16'b0000000011011000, 16'b1111111111110110, 16'b0000000000000000, 16'b1111111111101001, 16'b0000000000101001, 16'b1111111111101100, 16'b1111111111111111, 16'b0000000001010000, 16'b0000000001101100, 16'b1111111101110011, 16'b0000000001000111, 16'b0000000001011111, 16'b0000000000000110, 16'b0000000010101010, 16'b1111111110001100, 16'b1111111001100111, 16'b0000000000000000, 16'b1111111111111000, 16'b1111111111110010, 16'b1111111100000000, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111110011000, 16'b1111111111111000, 16'b1111111111001111, 16'b0000000001001111, 16'b0000000010111111, 16'b1111111111000010, 16'b1111111111100110, 16'b1111111111101011, 16'b0000000000001101, 16'b1111111100110111}, 
{16'b1111111110100101, 16'b0000000011000100, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000110010101, 16'b0000000010100100, 16'b1111111111111111, 16'b1111111011100011, 16'b0000000000111100, 16'b1111111010011010, 16'b1111110100110001, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000011011011, 16'b0000000000111000, 16'b0000000000000000, 16'b1111111101010111, 16'b0000000000000000, 16'b0000000000000011, 16'b0000000000011111, 16'b0000000001111100, 16'b1111111111110010, 16'b1111111101000111, 16'b0000000000000100, 16'b1111111111111010, 16'b0000001000101001, 16'b0000000010100111, 16'b1111111111111111, 16'b1111111111011011, 16'b0000000101010110, 16'b1111111111101011, 16'b1111111111010011}, 
{16'b1111111011110100, 16'b0000000001011001, 16'b1111111111101110, 16'b1111111111111111, 16'b1111111110000001, 16'b1111111100111110, 16'b0000000000011000, 16'b0000000001001001, 16'b1111111111111111, 16'b1111111110101000, 16'b1111111011011010, 16'b0000000001100110, 16'b0000000010011011, 16'b0000000000000000, 16'b0000000110101101, 16'b1111111011100000, 16'b0000000000110101, 16'b1111111100110111, 16'b0000000010010000, 16'b1111111111111111, 16'b1111111111101100, 16'b0000000000100011, 16'b0000000000111110, 16'b0000000000000000, 16'b1111111100000011, 16'b0000000000001111, 16'b1111111011100001, 16'b1111111111101011, 16'b1111111111111111, 16'b0000000101011001, 16'b1111111110011110, 16'b0000000000000000}, 
{16'b1111111111111111, 16'b0000000000111010, 16'b0000000000000000, 16'b0000000011001000, 16'b1111111111000100, 16'b1111111111101001, 16'b0000000000011101, 16'b1111111111111101, 16'b1111111111101000, 16'b0000000101001000, 16'b0000000101100101, 16'b0000000000000000, 16'b1111111101010101, 16'b1111111010011000, 16'b1111111111100110, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111011111, 16'b1111111100001100, 16'b0000000011000011, 16'b0000000000000001, 16'b0000000010111101, 16'b1111111111111111, 16'b0000000100011111, 16'b0000000000111111, 16'b0000000010011100, 16'b0000000011101001, 16'b1111111111100101, 16'b1111111100110111, 16'b1111111100011110, 16'b1111111111111101, 16'b1111111010101001}, 
{16'b1111111110001100, 16'b1111111111111111, 16'b0000000000111101, 16'b1111111100101001, 16'b0000000000101100, 16'b1111111111111111, 16'b1111111110010000, 16'b1111111111111011, 16'b1111111110111111, 16'b0000000000010011, 16'b0000000000100111, 16'b1111111111011011, 16'b0000000000001000, 16'b0000000001100000, 16'b1111111010111111, 16'b1111111110000010, 16'b0000000001110100, 16'b1111111110100101, 16'b0000000000000000, 16'b1111111111110011, 16'b0000000001100010, 16'b0000000000000100, 16'b1111111111110000, 16'b0000000000010101, 16'b0000000010001001, 16'b1111111111001010, 16'b0000000000000000, 16'b1111111100011000, 16'b1111111110011011, 16'b1111111111111100, 16'b0000000001011000, 16'b0000000000000000}, 
{16'b1111111011110101, 16'b0000000011010111, 16'b1111111111111111, 16'b1111111111111100, 16'b1111111111111011, 16'b0000000001011001, 16'b1111111111111111, 16'b0000000110001011, 16'b1111111111111000, 16'b1111111111111111, 16'b0000000001101001, 16'b0000000000010100, 16'b0000000000000011, 16'b0000000000000000, 16'b0000000000111110, 16'b0000000010101001, 16'b0000000001011011, 16'b0000000001010101, 16'b1111111111111011, 16'b0000000010011101, 16'b0000000000110011, 16'b0000000000010100, 16'b1111111111111011, 16'b0000000010000010, 16'b1111111111001101, 16'b1111111101010010, 16'b1111111111010000, 16'b1111111111111111, 16'b0000000000110100, 16'b0000000000001111, 16'b0000000001100100, 16'b0000000011110101}, 
{16'b1111111111110110, 16'b1111111100111000, 16'b0000000000011010, 16'b1111111111111111, 16'b0000000111010101, 16'b1111111110010101, 16'b1111111011011011, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111110010, 16'b0000000000011000, 16'b0000000011011111, 16'b0000000010100100, 16'b0000000000000101, 16'b0000000000010001, 16'b1111111110100110, 16'b0000000000010001, 16'b1111111111101100, 16'b0000000000000000, 16'b0000000000100110, 16'b1111111111101100, 16'b0000000000001001, 16'b0000000010001000, 16'b0000000000010010, 16'b1111111111111001, 16'b1111111100101100, 16'b0000000001101000, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111001001, 16'b1111111111110101, 16'b1111111111011111}, 
{16'b0000000000000011, 16'b1111111111011111, 16'b1111111110111111, 16'b1111111110010000, 16'b1111111011101000, 16'b0000000100111000, 16'b0000000000000000, 16'b0000000001010110, 16'b0000000010010010, 16'b0000000000000110, 16'b1111111111101110, 16'b0000000011110011, 16'b0000000001110010, 16'b1111111101000100, 16'b1111111110101100, 16'b1111111111101010, 16'b1111111100110100, 16'b1111111111110111, 16'b0000000000000000, 16'b1111111111111101, 16'b0000000001001111, 16'b1111111110111001, 16'b0000000000000000, 16'b0000000000100111, 16'b1111111111111111, 16'b1111111101010001, 16'b0000000001010000, 16'b0000000000000000, 16'b0000000000010110, 16'b0000000000000101, 16'b1111111101011110, 16'b0000000000001010}, 
{16'b1111111110011011, 16'b1111111110101111, 16'b0000000000100111, 16'b1111111111000000, 16'b1111111111010010, 16'b0000000000111011, 16'b1111111111111101, 16'b0000000000010001, 16'b0000000001000011, 16'b1111111111111111, 16'b0000000000111111, 16'b1111111110111110, 16'b1111111111111011, 16'b1111111111111111, 16'b0000000000110100, 16'b1111111111111111, 16'b0000000011111010, 16'b1111111111110111, 16'b0000000001111111, 16'b1111111110101001, 16'b0000000001010001, 16'b0000000000100000, 16'b0000000000101011, 16'b0000000000010010, 16'b1111111111010110, 16'b1111111101110001, 16'b1111111101111011, 16'b0000000000110111, 16'b1111111111010101, 16'b0000000000000000, 16'b1111111111110001, 16'b0000000001110110}, 
{16'b1111111111111111, 16'b1111111100110000, 16'b1111111100110100, 16'b1111111111111111, 16'b0000000101000011, 16'b1111111111010001, 16'b0000000000000000, 16'b0000000011110111, 16'b1111111110110100, 16'b0000000000000000, 16'b1111111100101010, 16'b1111111100000101, 16'b0000000011100101, 16'b0000000001001101, 16'b1111111111000001, 16'b1111111101110011, 16'b0000000001011000, 16'b0000000000000000, 16'b1111111110000110, 16'b0000000000001101, 16'b0000000000100011, 16'b1111111111010010, 16'b0000000010010001, 16'b1111111000001010, 16'b0000000000010100, 16'b0000000001111010, 16'b1111111111101010, 16'b0000000000000111, 16'b1111111110001000, 16'b1111111111111111, 16'b1111111110011001, 16'b1111111111110011}, 
{16'b0000000001101100, 16'b0000000010110000, 16'b0000000100011001, 16'b1111111110010111, 16'b0000000011010101, 16'b0000000010011100, 16'b0000000000000000, 16'b0000000011101001, 16'b0000000010110110, 16'b1111111111001001, 16'b0000000101100111, 16'b1111111101001101, 16'b0000000100111110, 16'b0000000011100100, 16'b1111110111011010, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000010, 16'b0000000010000101, 16'b1111111011111110, 16'b0000000001110001, 16'b1111111110010011, 16'b1111111100000100, 16'b1111111110101111, 16'b0000000010101000, 16'b1111111010101110, 16'b1111111101010111, 16'b1111111111101010, 16'b1111111111111111, 16'b1111111011011111, 16'b0000000011001010, 16'b0000000000000000}, 
{16'b1111111111100110, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111101001100, 16'b0000000000000100, 16'b0000000000000100, 16'b1111111111111000, 16'b1111111111110011, 16'b1111111111101000, 16'b0000000001000111, 16'b1111111111111111, 16'b0000000000101010, 16'b1111111101010000, 16'b0000000000110110, 16'b1111111111111111, 16'b0000000001001000, 16'b0000000011100101, 16'b1111111101001011, 16'b0000000000011010, 16'b1111111111001101, 16'b0000000001000001, 16'b0000000001100001, 16'b1111111111010100, 16'b1111111101111111, 16'b0000000000001010, 16'b0000000110101000, 16'b1111111111110011, 16'b1111111111111000, 16'b0000000010100110, 16'b0000000000000000, 16'b0000000110111001}, 
{16'b1111111011110100, 16'b0000000000010010, 16'b1111111110010001, 16'b0000000011000100, 16'b0000000000111000, 16'b1111111111101111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111101100100, 16'b1111111111101111, 16'b0000000000000000, 16'b1111111011100011, 16'b0000000000000110, 16'b1111111111101011, 16'b1111111111111110, 16'b1111111111111111, 16'b1111111111000100, 16'b0000000000000010, 16'b0000000000000001, 16'b0000000001010001, 16'b0000000000001000, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111011, 16'b0000000000000000, 16'b0000000000001001, 16'b0000000100101001, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111101011, 16'b0000000001011001, 16'b1111111111110010}, 
{16'b1111111111111111, 16'b1111111110110010, 16'b0000000001101000, 16'b0000000000010100, 16'b1111111101000001, 16'b0000000000000000, 16'b0000000010010010, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111001101, 16'b0000000000111010, 16'b0000000000001001, 16'b0000000010100101, 16'b1111111011100111, 16'b1111111111001111, 16'b1111111111110111, 16'b0000000001101110, 16'b1111111100111011, 16'b0000000000001010, 16'b1111111001111101, 16'b1111111111110110, 16'b1111111111000011, 16'b1111111111101011, 16'b0000000010010111, 16'b1111111111011001, 16'b1111111101110000, 16'b0000000000101110, 16'b0000000000000000, 16'b0000000011001010, 16'b0000000100001011, 16'b1111111101011000, 16'b1111111100011010}, 
{16'b0000000000100010, 16'b0000000000001101, 16'b1111111100101011, 16'b1111111111100010, 16'b1111111111111111, 16'b0000000000000001, 16'b0000000000110110, 16'b0000000011010010, 16'b0000000000000000, 16'b0000000000001010, 16'b0000000000100011, 16'b1111111011101011, 16'b1111111111011101, 16'b1111111011001010, 16'b0000000011110110, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111010110111, 16'b1111111111111111, 16'b1111111111011001, 16'b1111111111110101, 16'b0000000000000000, 16'b0000000000011111, 16'b1111111110110011, 16'b0000000000011011, 16'b0000000011010010, 16'b0000000011011010, 16'b0000000011000111, 16'b0000000010011101, 16'b0000000000000000, 16'b0000000000111010, 16'b0000000110010001}, 
{16'b1111111111110011, 16'b1111111110000110, 16'b0000000011000111, 16'b1111111111001011, 16'b0000000000100011, 16'b0000000001010101, 16'b1111111111111111, 16'b1111111101101101, 16'b1111111111010100, 16'b1111111011001100, 16'b0000000011100101, 16'b0000000000000001, 16'b0000000011010110, 16'b0000000101010111, 16'b1111111111000100, 16'b1111111001000010, 16'b1111111111001010, 16'b0000000011110000, 16'b1111111101101111, 16'b1111111110010101, 16'b0000000000011110, 16'b0000000000000000, 16'b1111111011101000, 16'b1111111110011110, 16'b1111111111101011, 16'b1111111111000001, 16'b0000000000111001, 16'b0000000101101000, 16'b0000000001111101, 16'b1111111111111111, 16'b0000000000101001, 16'b0000000000001110}, 
{16'b0000000000010101, 16'b0000000011101000, 16'b0000000000000000, 16'b0000000010010111, 16'b0000000110101001, 16'b1111111110101000, 16'b1111111111111111, 16'b1111111111101001, 16'b0000000010010110, 16'b1111111110011101, 16'b1111111111111111, 16'b0000000010101010, 16'b0000000000000100, 16'b0000000000001110, 16'b1111110011110010, 16'b1111111111010111, 16'b0000000000000000, 16'b0000000001100110, 16'b1111111111111110, 16'b0000000010011000, 16'b1111111111111111, 16'b1111111110100111, 16'b1111111011100000, 16'b0000000001000010, 16'b0000000010010010, 16'b1111110111001000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000100010110, 16'b1111111001100101, 16'b0000000000000000, 16'b1111111111111100}, 
{16'b0000000000000100, 16'b1111111101010010, 16'b0000000000011011, 16'b1111111111111000, 16'b0000000000011010, 16'b0000000100001110, 16'b1111111010001100, 16'b0000000000010001, 16'b0000000011011000, 16'b1111111101010011, 16'b1111111111110100, 16'b0000000000011001, 16'b1111111111111011, 16'b0000000001011011, 16'b0000000000110110, 16'b1111111111110111, 16'b0000000000100010, 16'b0000000000000000, 16'b0000000000001011, 16'b0000000011000010, 16'b1111111111110001, 16'b1111111100001000, 16'b1111111011001010, 16'b1111111110011100, 16'b1111111011010001, 16'b0000000001101010, 16'b0000000100111111, 16'b0000000010111100, 16'b1111111111111010, 16'b1111111101000001, 16'b1111111101100000, 16'b0000000000011110}, 
{16'b0000000000011010, 16'b1111111100001011, 16'b1111111111110111, 16'b0000000001001101, 16'b1111111100001011, 16'b0000000001010110, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000010000111, 16'b1111111111110111, 16'b0000000000000100, 16'b0000000000000000, 16'b0000000001000001, 16'b1111111111110111, 16'b0000000000000001, 16'b1111111111111111, 16'b1111111101011011, 16'b1111111011111101, 16'b1111111111111111, 16'b1111111011101110, 16'b1111111101100101, 16'b1111111101000001, 16'b0000000111000111, 16'b0000000000001001, 16'b1111111111101000, 16'b0000000010100010, 16'b0000000111001011, 16'b0000000011001010, 16'b1111110111100001, 16'b1111111110100001}, 
{16'b0000000011000000, 16'b1111111111111111, 16'b0000000010000000, 16'b1111111111110101, 16'b0000000011110111, 16'b1111111110110110, 16'b0000000000100100, 16'b0000000011010110, 16'b0000000010001001, 16'b1111111011110100, 16'b1111111111100000, 16'b0000000000111110, 16'b0000000000100011, 16'b1111111111111000, 16'b0000000000101011, 16'b0000000000000000, 16'b0000000010111001, 16'b0000000000010001, 16'b0000000010111111, 16'b1111111111011110, 16'b1111111110111110, 16'b1111111111011001, 16'b1111111111111111, 16'b0000000010011010, 16'b1111111110011000, 16'b1111111111111100, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000010010101, 16'b1111111101011011, 16'b1111111111110100}, 
{16'b1111111111111111, 16'b1111111111110000, 16'b1111111100010001, 16'b0000000010010001, 16'b0000000001110010, 16'b1111111111000111, 16'b1111111111111111, 16'b1111111110001011, 16'b0000000000000011, 16'b1111111111111111, 16'b1111111101100101, 16'b1111111110000001, 16'b0000000011110101, 16'b0000000000000000, 16'b1111111110111110, 16'b1111111111111111, 16'b0000000001101101, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111110010001, 16'b0000000010100001, 16'b0000000000000000, 16'b0000000001001111, 16'b1111111111110001, 16'b0000000001010000, 16'b0000000000000001, 16'b0000000000000000, 16'b0000000001111011, 16'b1111111110011101, 16'b1111111111101000, 16'b0000000001010010, 16'b1111111111001001}, 
{16'b1111111111110111, 16'b1111111101100010, 16'b0000000100110000, 16'b1111111111011110, 16'b0000000001100100, 16'b1111111101101101, 16'b0000000000000000, 16'b0000000000010001, 16'b1111111100001010, 16'b1111111111111001, 16'b1111111111000000, 16'b0000000000011101, 16'b1111111101011000, 16'b0000000001000110, 16'b0000000001100111, 16'b0000000000111000, 16'b0000000000101011, 16'b1111111111101100, 16'b1111111010010101, 16'b1111111111111001, 16'b1111111111100010, 16'b0000000001000111, 16'b1111111111000111, 16'b1111111111111111, 16'b0000000001100101, 16'b1111111111101000, 16'b1111111111111000, 16'b0000000011000111, 16'b1111111100110100, 16'b1111111101101000, 16'b0000000010110011, 16'b0000000000010010}, 
{16'b0000000011011100, 16'b0000000001100111, 16'b0000000000000000, 16'b1111111110101110, 16'b1111111111010111, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111011100, 16'b1111111111000000, 16'b1111111111000011, 16'b0000000000000000, 16'b0000000001010001, 16'b0000000000000011, 16'b0000000000011011, 16'b1111111111101001, 16'b0000000000000010, 16'b1111111110110001, 16'b0000000000000000, 16'b1111111111110110, 16'b1111111111111111, 16'b0000000000000001, 16'b0000000000011110, 16'b0000000000110001, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111011000111, 16'b1111111110011001, 16'b0000000000000011, 16'b0000000000001010, 16'b0000000000000000, 16'b1111111110100101, 16'b0000000000001010}, 
{16'b0000000001100000, 16'b1111110111101001, 16'b1111111111111111, 16'b1111111111011001, 16'b1111111110001000, 16'b1111111111111011, 16'b0000000000000000, 16'b0000000100011000, 16'b1111111111101001, 16'b1111111111110100, 16'b0000000000101010, 16'b1111111010101101, 16'b0000000000001100, 16'b1111111100011111, 16'b0000000101110001, 16'b1111111111100101, 16'b1111111110001100, 16'b1111111011100111, 16'b1111111111111010, 16'b1111111010010101, 16'b1111111001100001, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000001111100, 16'b1111111111111000, 16'b1111111101100111, 16'b1111111111011010, 16'b1111111111110100, 16'b0000000000000000, 16'b1111111111101111, 16'b1111111010011001}
};

localparam logic signed [15:0] bias [32] = '{
16'b0000000010000111,  // 0.5280959606170654
16'b0000000011010111,  // 0.8414360880851746
16'b0000000001100101,  // 0.397830605506897
16'b0000000001101001,  // 0.4105983078479767
16'b1111110001010111,  // -3.657735586166382
16'b1111111100011010,  // -0.8977976441383362
16'b0000000110110100,  // 1.7051936388015747
16'b1111111010111001,  // -1.2765135765075684
16'b1111111101101010,  // -0.5837795734405518
16'b0000001010110011,  // 2.699671983718872
16'b0000000000110111,  // 0.2170683741569519
16'b0000000011100001,  // 0.8814588785171509
16'b1111110101011101,  // -2.634300947189331
16'b1111111000011111,  // -1.877297282218933
16'b0000000110101001,  // 1.6625694036483765
16'b0000001010111110,  // 2.7459704875946045
16'b1111111110000101,  // -0.47838035225868225
16'b0000000110110010,  // 1.6984987258911133
16'b0000000011011010,  // 0.8548859357833862
16'b0000000100000001,  // 1.0045719146728516
16'b0000000101101011,  // 1.4197649955749512
16'b0000000011010101,  // 0.832463800907135
16'b0000000010001011,  // 0.5434179306030273
16'b0000000011101101,  // 0.9277304410934448
16'b1111111110101000,  // -0.3426123857498169
16'b1111111101110000,  // -0.5587119460105896
16'b1111111101100001,  // -0.6208624839782715
16'b1111111010111000,  // -1.2802538871765137
16'b0000000000001111,  // 0.05940237268805504
16'b1111111100101101,  // -0.8213341236114502
16'b0000000011100000,  // 0.8783953189849854
16'b1111111100001100   // -0.949700653553009
};
endpackage