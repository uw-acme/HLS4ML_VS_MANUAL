// Package with weights and biases for reset gate dense latency layer
`ifndef RESET_GATE_PKG
    `define RESET_GATE_PKG reset_gate
`endif

// Package with weights and biases for update gate dense latency layer
`ifndef UPDATE_GATE_PKG
    `define UPDATE_GATE_PKG update_gate
`endif

// Package with weights and biases for candidate gate dense latency layer
`ifndef CANDIDATE_HIDDEN_STATE_PKG
    `define CANDIDATE_HIDDEN_STATE_PKG candidate_hidden_state
`endif
