// Width: 28
// NFRAC: 14
package dense_1_28_14;

localparam logic signed [27:0] weights [16][64] = '{ 
{28'b0000000000000001000001010010, 28'b1111111111111101011001001001, 28'b1111111111111111010001101111, 28'b1111111111111111000110000001, 28'b1111111111111110011000010100, 28'b0000000000000000011100010000, 28'b1111111111111011110110100001, 28'b0000000000000000000000000001, 28'b0000000000000000001110110111, 28'b0000000000000001000011011101, 28'b0000000000000000000000110000, 28'b1111111111111110011000011011, 28'b1111111111111111111111101110, 28'b0000000000000000110101100001, 28'b0000000000000000001000100100, 28'b1111111111111110111101000001, 28'b0000000000000000111011100110, 28'b0000000000000000001111000001, 28'b0000000000000000000000000001, 28'b1111111111111111111111111101, 28'b0000000000000001100000011111, 28'b1111111111111110101011001001, 28'b1111111111111111111010010110, 28'b0000000000000001111001000000, 28'b1111111111111110101101101100, 28'b1111111111111101010001010000, 28'b1111111111111110111001011111, 28'b1111111111111111001110000001, 28'b1111111111111111100101001110, 28'b1111111111111111111111100011, 28'b0000000000000000001001101010, 28'b0000000000000000111110110100, 28'b0000000000000000110010000111, 28'b1111111111111111111100101001, 28'b0000000000000000000000000010, 28'b0000000000000001001111101110, 28'b1111111111111111111011011000, 28'b1111111111111110111111101100, 28'b0000000000000000000110111110, 28'b0000000000000000110001010010, 28'b1111111111111111111100111011, 28'b0000000000000001000110011100, 28'b1111111111111110111011110011, 28'b0000000000000011101101110000, 28'b1111111111111111111111101110, 28'b0000000000000001110011110110, 28'b0000000000000000000000000000, 28'b0000000000000000101111001100, 28'b0000000000000000110010001100, 28'b1111111111111111111001111111, 28'b0000000000000000000000000000, 28'b0000000000000000101001000100, 28'b0000000000000000110111010001, 28'b0000000000000000010011111010, 28'b1111111111111111100010011111, 28'b1111111111111110110000100011, 28'b0000000000000010001001010100, 28'b1111111111111110000000000110, 28'b0000000000000001110111101110, 28'b1111111111111110100101010010, 28'b0000000000000011001011000010, 28'b1111111111111111111110000111, 28'b0000000000000000000010111011, 28'b0000000000000000010100110001}, 
{28'b0000000000000000000000101110, 28'b1111111111111110101101111000, 28'b1111111111111111011110000110, 28'b1111111111111110111000011011, 28'b1111111111111110101110101111, 28'b0000000000000000011011010011, 28'b1111111111111100111110110111, 28'b1111111111111111111111011011, 28'b1111111111111111000101110100, 28'b0000000000000000101100001000, 28'b0000000000000000000001101100, 28'b1111111111111111101001111100, 28'b0000000000000000110010011101, 28'b0000000000000000000000000001, 28'b1111111111111111111111111101, 28'b0000000000000000110101001001, 28'b1111111111111111111110011101, 28'b0000000000000000000000000101, 28'b1111111111111111010001010111, 28'b1111111111111110111111111100, 28'b0000000000000001110001001111, 28'b1111111111111111101011010010, 28'b0000000000000000001100010001, 28'b0000000000000010110010111010, 28'b0000000000000001000001111011, 28'b1111111111111111000101000010, 28'b1111111111111111000100111000, 28'b1111111111111111111111111010, 28'b1111111111111111100110000001, 28'b1111111111111110011000001111, 28'b1111111111111111110000101011, 28'b0000000000000001110100011101, 28'b0000000000000001000111010100, 28'b0000000000000010001100110101, 28'b0000000000000010100001000010, 28'b0000000000000000001100111011, 28'b1111111111111111100001101100, 28'b1111111111111110010000111001, 28'b0000000000000000001110100000, 28'b0000000000000000110000010110, 28'b0000000000000000000101110111, 28'b0000000000000000110100110110, 28'b1111111111111111001001100100, 28'b0000000000000001000000100000, 28'b0000000000000000101100000111, 28'b0000000000000000001100110000, 28'b1111111111111110101000111110, 28'b0000000000000000010100010110, 28'b0000000000000001000010101111, 28'b0000000000000000000111101010, 28'b0000000000000000000110010111, 28'b0000000000000100101000010000, 28'b1111111111111111101100110111, 28'b1111111111111111100110111010, 28'b1111111111111111110010000110, 28'b1111111111111111111110000000, 28'b0000000000000001000001110001, 28'b1111111111111110100001010011, 28'b0000000000000011111100001111, 28'b0000000000000000000001001110, 28'b0000000000000010000101010001, 28'b0000000000000000111101011111, 28'b0000000000000011010010100111, 28'b0000000000000000100100000110}, 
{28'b1111111111111111111110000011, 28'b0000000000000000000000000000, 28'b1111111111111111101010101101, 28'b1111111111111111010010111100, 28'b1111111111111111010000101111, 28'b0000000000000000001010101101, 28'b0000000000000101111011000111, 28'b1111111111111111111111111111, 28'b1111111111111010111011111001, 28'b1111111111111111111111111110, 28'b1111111111111111111111100011, 28'b1111111111111111111011011010, 28'b1111111111111111000101110010, 28'b0000000000000000000000010100, 28'b1111111111111111111101100110, 28'b0000000000000000101011000010, 28'b0000000000000011100111110010, 28'b1111111111111111111111111111, 28'b0000000000000000010010011111, 28'b0000000000000000000000000101, 28'b0000000000000001101001100001, 28'b1111111111111101000111010111, 28'b0000000000000010010011110101, 28'b1111111111111101001001010010, 28'b0000000000000011110010110100, 28'b1111111111111110100111010100, 28'b1111111111111111000001010101, 28'b1111111111111101001000010011, 28'b0000000000000101000110000001, 28'b0000000000000001000110100111, 28'b0000000000000000000010111010, 28'b0000000000000010000100100010, 28'b0000000000000100000101001110, 28'b1111111111111011001110000101, 28'b1111111111111111100111100010, 28'b0000000000000000001000001011, 28'b1111111111111111000100110111, 28'b0000000000000011100101101000, 28'b1111111111111111110101111011, 28'b0000000000000001010000001001, 28'b0000000000000001010101010001, 28'b0000000000000001011110101001, 28'b1111111111111111111111111111, 28'b1111111111111111111111111101, 28'b1111111111111111111011100101, 28'b0000000000000000101000001110, 28'b1111111111111110111000011000, 28'b1111111111111111010100011010, 28'b1111111111111111111011100010, 28'b0000000000000001100100101100, 28'b1111111111111111010010111101, 28'b0000000000000000100110011100, 28'b1111111111111111111111111000, 28'b0000000000000000100010010111, 28'b1111111111111111010011000100, 28'b1111111111111111111111111110, 28'b1111111111111110110001000100, 28'b1111111111111101010100100110, 28'b1111111111111111111111011111, 28'b0000000000000000000000000000, 28'b0000000000000110001010111110, 28'b0000000000000000000011010101, 28'b1111111111111111111111010100, 28'b1111111111111110110000110010}, 
{28'b1111111111111110001010101101, 28'b1111111111111110100001101001, 28'b1111111111111101001110101011, 28'b0000000000000001001110111010, 28'b1111111111111110101111001000, 28'b1111111111111010100111010111, 28'b1111111111111111100010101000, 28'b1111111111111110110001001000, 28'b0000000000000000111001010111, 28'b1111111111111111111111111111, 28'b0000000000000101000011111100, 28'b1111111111111111100100111111, 28'b1111111111111100110111101100, 28'b0000000000000010010100010010, 28'b0000000000000000000110011100, 28'b1111111111111111111111100111, 28'b1111111111111110001110011001, 28'b1111111111111111111111111111, 28'b0000000000000000000000000001, 28'b1111111111111111000110000111, 28'b1111111111111011011001010111, 28'b1111111111111111100011011011, 28'b1111111111111101001101001111, 28'b0000000000000000110010110011, 28'b1111111111111110011100111110, 28'b1111111111111100010100010100, 28'b0000000000000001010000000100, 28'b0000000000000010111100100100, 28'b0000000000000101001011100101, 28'b1111111111111110001010010000, 28'b1111111111111101101010110110, 28'b0000000000000000010010111010, 28'b0000000000000010000000000010, 28'b1111111111111100101000101000, 28'b1111111111111110101111100000, 28'b0000000000000000000000000000, 28'b1111111111111101000110001000, 28'b0000000000000000111110000101, 28'b1111111111111110001111000100, 28'b0000000000000000011110100011, 28'b0000000000000001110101011001, 28'b0000000000000000101000001000, 28'b0000000000000000000000000000, 28'b0000000000000000000101001101, 28'b0000000000000010001101011100, 28'b1111111111111111001100110100, 28'b1111111111111111111111111110, 28'b1111111111111110100111111100, 28'b1111111111111111111111111110, 28'b1111111111111111100111001111, 28'b1111111111111101100010011101, 28'b0000000000000000010110001110, 28'b1111111111111111111111111110, 28'b0000000000000000110111110110, 28'b0000000000000001010000101111, 28'b0000000000000010100101101010, 28'b1111111111111100001000010011, 28'b1111111111111100010010001110, 28'b1111111111111101001011011111, 28'b0000000000000011011101110000, 28'b0000000000000110111111110001, 28'b1111111111111100011001101100, 28'b1111111111111111110010001001, 28'b0000000000000001101111001011}, 
{28'b0000000000000001010111100110, 28'b1111111111111101100001101011, 28'b1111111111111110111101100111, 28'b1111111111111111111111111111, 28'b1111111111111111011000100101, 28'b0000000000000001010111000110, 28'b0000000000000000110000100000, 28'b1111111111111111111111111101, 28'b1111111111111101100111000101, 28'b1111111111111111000010000111, 28'b1111111111111110100001100111, 28'b0000000000000000001101100011, 28'b0000000000000000000000010100, 28'b0000000000000000000000000000, 28'b1111111111111111110101101000, 28'b0000000000000001011011100011, 28'b0000000000000000100010001101, 28'b1111111111111110011011011011, 28'b0000000000000000000111110110, 28'b0000000000000000000011011101, 28'b0000000000000000110101110011, 28'b1111111111111111100001110010, 28'b0000000000000000010011000011, 28'b1111111111111111111011000111, 28'b0000000000000100010000110110, 28'b1111111111111111010000010011, 28'b1111111111111110111000000001, 28'b1111111111111110011000101010, 28'b0000000000000000000000000001, 28'b0000000000000000101010001011, 28'b0000000000000000011101110000, 28'b0000000000000001000110000010, 28'b1111111111111111111100110100, 28'b0000000000000000010010111110, 28'b0000000000000000100001011101, 28'b1111111111111111111111111111, 28'b0000000000000000000001100101, 28'b0000000000000011100001101011, 28'b1111111111111110110110000011, 28'b1111111111111111101100011000, 28'b0000000000000001101110111010, 28'b0000000000000000111111101100, 28'b1111111111111110000010110101, 28'b0000000000000000000001100000, 28'b1111111111111011101110100000, 28'b1111111111111111111111111111, 28'b1111111111111111100000101000, 28'b0000000000000000000011000011, 28'b1111111111111111111111111101, 28'b1111111111111111111001111111, 28'b1111111111111111111111111111, 28'b0000000000000000110000001001, 28'b1111111111111111111110101100, 28'b0000000000000001010001010110, 28'b1111111111111111001111000100, 28'b1111111111111101000011110011, 28'b1111111111111110001000100110, 28'b1111111111111101111101100110, 28'b1111111111111101100010110110, 28'b0000000000000010111111001101, 28'b0000000000000101011111101001, 28'b0000000000000011001010111110, 28'b0000000000000000011111011000, 28'b1111111111111111111111111101}, 
{28'b1111111111111110001101111011, 28'b1111111111111101011110100100, 28'b0000000000000000000000000010, 28'b0000000000000001001110101001, 28'b0000000000000001001001000010, 28'b1111111111111111001001101101, 28'b0000000000000010010101000010, 28'b1111111111111111111111111110, 28'b0000000000000000111110011000, 28'b1111111111111111111111111111, 28'b1111111111111111111101100110, 28'b1111111111111111101101011010, 28'b1111111111111111010010110101, 28'b0000000000000010010100000000, 28'b1111111111111111101001001001, 28'b0000000000000000000000000011, 28'b1111111111111101100000000010, 28'b1111111111111110100101010001, 28'b0000000000000000000000000010, 28'b1111111111111111111111111110, 28'b1111111111111111110011110100, 28'b1111111111111110101111101010, 28'b1111111111111110101110011001, 28'b0000000000000001110111001001, 28'b1111111111111110101110100101, 28'b1111111111111111111111110001, 28'b0000000000000001000001100100, 28'b1111111111111111101101010011, 28'b1111111111111100010001001101, 28'b1111111111111111111111111110, 28'b1111111111111111101110111000, 28'b1111111111111111111101010111, 28'b1111111111111111111101000010, 28'b0000000000000000001010011110, 28'b0000000000000000100001110001, 28'b0000000000000001011000100000, 28'b0000000000000000000011011110, 28'b1111111111111111100110111001, 28'b1111111111111110111100110001, 28'b1111111111111111111111100001, 28'b1111111111111111010100101110, 28'b1111111111111101111001111001, 28'b0000000000000001100110011111, 28'b0000000000000000000010110000, 28'b0000000000000010011010011101, 28'b0000000000000000000000000000, 28'b1111111111111111111111111101, 28'b0000000000000000011000010101, 28'b1111111111111110010100101100, 28'b0000000000000000111011111010, 28'b0000000000000000000000000000, 28'b1111111111111111100110001000, 28'b1111111111111110100011011111, 28'b0000000000000001100010111100, 28'b1111111111111111111111111111, 28'b0000000000000001011000110110, 28'b0000000000000000110111011101, 28'b0000000000000000110100001100, 28'b1111111111111111111011001110, 28'b1111111111111111111101111000, 28'b1111111111111100110001000101, 28'b1111111111111111011111101100, 28'b1111111111111111110001011000, 28'b1111111111111111111111111001}, 
{28'b1111111111111110110111100110, 28'b1111111111111110101010001101, 28'b1111111111111110010001100001, 28'b1111111111111111101110001100, 28'b1111111111111111011101111000, 28'b0000000000000000011010101100, 28'b1111111111111101001101010001, 28'b1111111111111111011001100101, 28'b1111111111111111000110100101, 28'b1111111111111111111111111101, 28'b1111111111111110110110011010, 28'b0000000000000001011001000100, 28'b0000000000000000001001000111, 28'b0000000000000000100011010001, 28'b0000000000000001001111110111, 28'b0000000000000000000000000100, 28'b0000000000000011001100000101, 28'b0000000000000000010110111000, 28'b0000000000000000111110001010, 28'b0000000000000001000100101110, 28'b1111111111111111010111111000, 28'b0000000000000001011101000001, 28'b1111111111111111000001111000, 28'b1111111111111101111111100000, 28'b0000000000000000101100011000, 28'b0000000000000010000100010010, 28'b1111111111111111111110111011, 28'b0000000000000000001101110010, 28'b1111111111111100001100100101, 28'b0000000000000001001001010110, 28'b0000000000000001000100011001, 28'b1111111111111110100000011100, 28'b0000000000000001111000101100, 28'b0000000000000010101010001010, 28'b0000000000000000000000000000, 28'b0000000000000001010111101001, 28'b1111111111111111111111111111, 28'b0000000000000001001000110001, 28'b0000000000000000110010111110, 28'b0000000000000000000000000000, 28'b1111111111111111100001110100, 28'b1111111111111110100010111010, 28'b0000000000000000100100101110, 28'b0000000000000001111011101111, 28'b0000000000000010000100111000, 28'b1111111111111111010100111101, 28'b1111111111111111101010101000, 28'b1111111111111111001111011001, 28'b1111111111111111011101011000, 28'b0000000000000000011110010011, 28'b0000000000000000000000110100, 28'b0000000000000000001000101110, 28'b0000000000000000000000000000, 28'b0000000000000000101110011011, 28'b1111111111111111010011010100, 28'b0000000000000011000101010110, 28'b0000000000000001011011001000, 28'b1111111111111111111001101011, 28'b0000000000000001100011111010, 28'b0000000000000000110111100100, 28'b1111111111111001011111111111, 28'b1111111111111101101100011110, 28'b1111111111111111010011111010, 28'b1111111111111111111101011100}, 
{28'b0000000000000000000001010100, 28'b0000000000000000111101001111, 28'b1111111111111111111111111010, 28'b1111111111111111111111110111, 28'b1111111111111110101101100001, 28'b1111111111111111111000000000, 28'b1111111111111110111110000111, 28'b0000000000000000000000000001, 28'b0000000000000000000111000011, 28'b0000000000000001100011100010, 28'b0000000000000000000011101111, 28'b1111111111111110011111010000, 28'b1111111111111111101111111111, 28'b0000000000000000000000000010, 28'b1111111111111111110010100000, 28'b1111111111111110001100111001, 28'b1111111111111100100110110011, 28'b1111111111111111111111111011, 28'b1111111111111101100101010011, 28'b1111111111111110001101110110, 28'b1111111111111110011100010010, 28'b0000000000000001011000111000, 28'b0000000000000000001100000001, 28'b1111111111111111011011100010, 28'b1111111111111110010000001000, 28'b0000000000000000100111110010, 28'b0000000000000000000000000000, 28'b0000000000000001111111110101, 28'b0000000000000011001110010101, 28'b1111111111111111110101101101, 28'b0000000000000000000000001011, 28'b0000000000000000111011000001, 28'b1111111111111101010001010111, 28'b1111111111111110100001000011, 28'b0000000000000000001110001110, 28'b0000000000000000010111101101, 28'b1111111111111110111000001011, 28'b0000000000000000111101010100, 28'b0000000000000000100001110011, 28'b1111111111111111011000111001, 28'b1111111111111110010100100001, 28'b1111111111111111110110100001, 28'b0000000000000000001000011001, 28'b1111111111111111010101011110, 28'b0000000000000000001110010010, 28'b0000000000000000111010101101, 28'b1111111111111111100001011100, 28'b0000000000000000000110000111, 28'b0000000000000000000000000000, 28'b1111111111111111001000001111, 28'b1111111111111110011100100111, 28'b0000000000000001101010011111, 28'b0000000000000000100000011111, 28'b1111111111111111010010011001, 28'b0000000000000000100001111011, 28'b1111111111111111110000001101, 28'b1111111111111110000110100010, 28'b1111111111111111011101111000, 28'b1111111111111111110010101000, 28'b1111111111111111101110000010, 28'b0000000000000011010100100101, 28'b0000000000000000110000110111, 28'b1111111111111111110011100110, 28'b1111111111111111111111111010}, 
{28'b0000000000000000000011110000, 28'b0000000000000010010110001111, 28'b1111111111111101101011010110, 28'b1111111111111111000100110110, 28'b0000000000000001010010100110, 28'b1111111111111111001011001111, 28'b0000000000000100110110000100, 28'b1111111111111110110110010110, 28'b1111111111111111111111111101, 28'b0000000000000001001011000100, 28'b0000000000000001000001000101, 28'b1111111111111111111111010111, 28'b1111111111111111110011101101, 28'b1111111111111110000100100101, 28'b0000000000000001001000000010, 28'b0000000000000000101000111001, 28'b1111111111111111001110011000, 28'b1111111111111111111111111111, 28'b0000000000000000000000000000, 28'b0000000000000000000000000100, 28'b0000000000000001000011111011, 28'b1111111111111110001010010100, 28'b0000000000000001100100011001, 28'b0000000000000010011100111000, 28'b1111111111111111101001101010, 28'b1111111111111111111111111011, 28'b1111111111111111111011110101, 28'b1111111111111111111111111100, 28'b0000000000000010111100011101, 28'b0000000000000000000001010001, 28'b1111111111111110111010000011, 28'b0000000000000000000000000000, 28'b0000000000000001100010010110, 28'b1111111111111100110000011000, 28'b1111111111111101110101100101, 28'b0000000000000000110010111000, 28'b0000000000000000100011011101, 28'b1111111111111101101101101101, 28'b1111111111111111001111100100, 28'b1111111111111111001001001010, 28'b0000000000000001100110101010, 28'b0000000000000001100100000101, 28'b0000000000000000000000000001, 28'b1111111111111110111010111000, 28'b0000000000000000000000001101, 28'b0000000000000001100101001110, 28'b1111111111111111110000111010, 28'b1111111111111111111111111101, 28'b0000000000000000000010111100, 28'b0000000000000000111110101110, 28'b1111111111111111110001010011, 28'b1111111111111111001110011100, 28'b0000000000000001011000000111, 28'b1111111111111111001000111101, 28'b0000000000000001000111100110, 28'b0000000000000010010101101011, 28'b0000000000000000001010001111, 28'b0000000000000001000011011110, 28'b1111111111111110011001100011, 28'b1111111111111110100010000100, 28'b0000000000000011010100111101, 28'b1111111111111111011111000010, 28'b0000000000000000001011110000, 28'b1111111111111111101000000100}, 
{28'b0000000000000000000100001001, 28'b1111111111111110001100001011, 28'b0000000000000001011110011011, 28'b1111111111111110110111010100, 28'b1111111111111111111111001111, 28'b0000000000000000110110001001, 28'b1111111111111101101011000001, 28'b0000000000000000110001000000, 28'b0000000000000001111101100100, 28'b0000000000000000100111011110, 28'b0000000000000001011100110000, 28'b0000000000000001010010100100, 28'b1111111111111110110001111111, 28'b1111111111111111101100100100, 28'b1111111111111111110010110101, 28'b0000000000000000000000010011, 28'b1111111111111100001010010100, 28'b0000000000000001010010101110, 28'b1111111111111111110110101111, 28'b0000000000000000000111111101, 28'b1111111111111110100101110000, 28'b0000000000000000010001111000, 28'b0000000000000000100111001100, 28'b1111111111111111111111111010, 28'b1111111111111110001010001011, 28'b1111111111111111110011110001, 28'b1111111111111111101011000000, 28'b0000000000000100111111011101, 28'b1111111111111101010110011001, 28'b0000000000000000010001000000, 28'b0000000000000000011000110101, 28'b1111111111111111110001000010, 28'b1111111111111111000111011100, 28'b0000000000000000011101110101, 28'b1111111111111111101011111110, 28'b1111111111111111011101100110, 28'b1111111111111111010010011011, 28'b1111111111111111001010001110, 28'b1111111111111111111010010110, 28'b1111111111111110110011110110, 28'b0000000000000001010010011000, 28'b0000000000000000011111100110, 28'b0000000000000001111111001011, 28'b0000000000000000010110011101, 28'b0000000000000000001001011100, 28'b1111111111111110110101100010, 28'b0000000000000000000000000000, 28'b1111111111111111111111111101, 28'b1111111111111111111111111000, 28'b0000000000000000110001100111, 28'b0000000000000000101101011011, 28'b0000000000000001001011011111, 28'b1111111111111111111110011100, 28'b1111111111111110110100111001, 28'b0000000000000000000010010011, 28'b0000000000000000000000000001, 28'b0000000000000001010010100011, 28'b1111111111111111001100100100, 28'b1111111111111101110011000101, 28'b0000000000000010001111101100, 28'b1111111111111110110100110001, 28'b0000000000000100101001111100, 28'b1111111111111111111010111011, 28'b1111111111111110100101010000}, 
{28'b1111111111111101101100011111, 28'b1111111111111111111111100001, 28'b1111111111111110010111001001, 28'b0000000000000000111010111111, 28'b0000000000000001000011011011, 28'b1111111111111111100101110011, 28'b0000000000000010000100010110, 28'b1111111111111111010100011000, 28'b1111111111111110000101010010, 28'b1111111111111110100010000100, 28'b1111111111111110111111101100, 28'b1111111111111110000110001011, 28'b1111111111111111000101011001, 28'b0000000000000000110010011010, 28'b0000000000000000000000000000, 28'b0000000000000000000000000100, 28'b0000000000000011010111101100, 28'b1111111111111111110100111100, 28'b1111111111111111111111101110, 28'b0000000000000001101001010001, 28'b0000000000000001001010111101, 28'b1111111111111101101011110111, 28'b1111111111111110011110000111, 28'b0000000000000000110000011001, 28'b1111111111111110010001110001, 28'b1111111111111111111010101000, 28'b1111111111111110111101100011, 28'b1111111111111110101010011101, 28'b1111111111111110010000011110, 28'b0000000000000001001101010111, 28'b0000000000000000111010010100, 28'b1111111111111111011000000101, 28'b1111111111111111101101011001, 28'b1111111111111100000110101010, 28'b1111111111111111010010110001, 28'b0000000000000000001100101010, 28'b1111111111111111011110110101, 28'b1111111111111110110100000110, 28'b1111111111111111111111000100, 28'b0000000000000000011110011100, 28'b1111111111111111100001100000, 28'b1111111111111111111111010101, 28'b1111111111111111110111000011, 28'b1111111111111101010101111111, 28'b0000000000000000000000001101, 28'b0000000000000000000000000000, 28'b0000000000000001010111000100, 28'b1111111111111111100000001011, 28'b0000000000000001101100011101, 28'b1111111111111111001111001110, 28'b0000000000000001001001101111, 28'b1111111111111111111111101000, 28'b0000000000000000111001110011, 28'b1111111111111110011011110101, 28'b1111111111111111111111111111, 28'b0000000000000010000011000100, 28'b0000000000000001010000000011, 28'b0000000000000001001010110001, 28'b0000000000000000000110011111, 28'b1111111111111110011001101001, 28'b1111111111111110110011011101, 28'b1111111111111101010000010111, 28'b1111111111111111111111100001, 28'b0000000000000000011011011011}, 
{28'b0000000000000001001110111110, 28'b0000000000000000000000101010, 28'b0000000000000000100001100100, 28'b1111111111111111111111111111, 28'b0000000000000000100111010010, 28'b1111111111111111011101100000, 28'b0000000000000000111100000111, 28'b0000000000000000001010110111, 28'b0000000000000000100010110001, 28'b0000000000000001010111000011, 28'b1111111111111110111100100011, 28'b1111111111111111111010101100, 28'b1111111111111111111101111000, 28'b1111111111111111111101110000, 28'b1111111111111101010111000101, 28'b1111111111111110110011110001, 28'b0000000000000010100001011011, 28'b1111111111111111111000110110, 28'b1111111111111111110010101010, 28'b0000000000000000000000000100, 28'b1111111111111110011110101011, 28'b0000000000000000000010010101, 28'b0000000000000001000000001111, 28'b0000000000000000001001101111, 28'b0000000000000000001001011010, 28'b0000000000000001010110101000, 28'b0000000000000000000000000000, 28'b0000000000000000001001101000, 28'b0000000000000000000000000000, 28'b1111111111111111110011111000, 28'b1111111111111111001100100111, 28'b1111111111111101010101100010, 28'b0000000000000001000011101000, 28'b0000000000000001010111110011, 28'b1111111111111111111000100000, 28'b1111111111111111000011111011, 28'b0000000000000000000000000000, 28'b1111111111111101011000011010, 28'b1111111111111111110100010010, 28'b1111111111111111111111001011, 28'b0000000000000000110010001011, 28'b1111111111111111011110100101, 28'b1111111111111111111111111110, 28'b0000000000000011011000111011, 28'b0000000000000001110010110000, 28'b1111111111111111111110011111, 28'b1111111111111111111111111010, 28'b1111111111111111111111111110, 28'b1111111111111111000010011011, 28'b0000000000000000100101101001, 28'b0000000000000000100100111000, 28'b0000000000000000101100101110, 28'b0000000000000000101000010010, 28'b0000000000000001100011011001, 28'b0000000000000001011001100010, 28'b0000000000000010101000110100, 28'b1111111111111111011100001101, 28'b0000000000000001100100101100, 28'b0000000000000000100111000110, 28'b1111111111111110101100100111, 28'b0000000000000000011100011000, 28'b1111111111111110011100100100, 28'b1111111111111110001111011011, 28'b1111111111111110000000010110}, 
{28'b0000000000000000000000000101, 28'b0000000000000000111010011110, 28'b1111111111111111001110001011, 28'b0000000000000000000000000001, 28'b1111111111111111110011011100, 28'b1111111111111111110111010001, 28'b1111111111111101010110111010, 28'b1111111111111111111111111110, 28'b0000000000000001000000111000, 28'b0000000000000000111111111101, 28'b0000000000000000111100110111, 28'b1111111111111110011010000101, 28'b1111111111111111101001001010, 28'b0000000000000001001000101101, 28'b1111111111111111111111111011, 28'b0000000000000000000001001110, 28'b1111111111111100101000100110, 28'b1111111111111111111111111010, 28'b0000000000000001011111010111, 28'b0000000000000000010010000011, 28'b0000000000000000111100111101, 28'b1111111111111111100010011111, 28'b0000000000000000111111111010, 28'b0000000000000001100111101010, 28'b1111111111111110100101000011, 28'b1111111111111110111000011001, 28'b1111111111111111111110101100, 28'b1111111111111111101011010100, 28'b0000000000000000010001001101, 28'b0000000000000000000000000010, 28'b1111111111111111111111111110, 28'b0000000000000001010000011100, 28'b1111111111111101000000000011, 28'b0000000000000001011100100000, 28'b0000000000000010000000010111, 28'b0000000000000000011101110101, 28'b0000000000000000011100110010, 28'b1111111111111111100100010111, 28'b0000000000000000011101011111, 28'b1111111111111111100100101011, 28'b1111111111111110111111101100, 28'b1111111111111111110011000111, 28'b0000000000000000101010000110, 28'b0000000000000010110011000010, 28'b1111111111111100100111000011, 28'b1111111111111110001101111001, 28'b0000000000000000110001001011, 28'b1111111111111111100110111100, 28'b0000000000000001110011010110, 28'b1111111111111111000011100011, 28'b1111111111111110101011010000, 28'b1111111111111110111000010000, 28'b1111111111111111111111111111, 28'b0000000000000000011110110010, 28'b1111111111111111010111101111, 28'b1111111111111100101001110100, 28'b1111111111111111011011011001, 28'b1111111111111111111101011000, 28'b0000000000000000001011001001, 28'b1111111111111101100011110001, 28'b0000000000000100011110101111, 28'b1111111111111101110100101010, 28'b0000000000000010001010101011, 28'b0000000000000000100111001110}, 
{28'b0000000000000000010100000010, 28'b1111111111111111001110111010, 28'b0000000000000010100000110100, 28'b1111111111111110110010100111, 28'b1111111111111110001001011000, 28'b0000000000000000010111000000, 28'b0000000000000001001111001101, 28'b0000000000000001001100111110, 28'b1111111111111111010010100100, 28'b1111111111111111010110111001, 28'b0000000000000000001101011100, 28'b0000000000000000111010101001, 28'b0000000000000000111100001000, 28'b0000000000000000001100110110, 28'b1111111111111111001011101110, 28'b0000000000000000100000111000, 28'b0000000000000001111000100000, 28'b1111111111111111111101001001, 28'b1111111111111110111000011001, 28'b0000000000000000000000000010, 28'b0000000000000000010011000011, 28'b0000000000000000000101001100, 28'b1111111111111110110100111101, 28'b0000000000000000011100111010, 28'b0000000000000011001001011111, 28'b0000000000000000000010100100, 28'b0000000000000000101110001111, 28'b1111111111111100110100111101, 28'b1111111111111111101101011001, 28'b0000000000000000000010011000, 28'b1111111111111111001101110001, 28'b1111111111111110110000001110, 28'b0000000000000001110101010100, 28'b1111111111111111111001001100, 28'b1111111111111111110110010110, 28'b1111111111111110110001111001, 28'b0000000000000000100011011100, 28'b0000000000000001001010110010, 28'b1111111111111111111101100010, 28'b1111111111111111110100111000, 28'b1111111111111111010000001110, 28'b0000000000000000111010011100, 28'b0000000000000000000000000001, 28'b1111111111111101010000010011, 28'b0000000000000001001111101011, 28'b0000000000000001100110001001, 28'b1111111111111111111111111100, 28'b0000000000000000000110100001, 28'b1111111111111110010000111011, 28'b1111111111111111101100110100, 28'b1111111111111111111111111111, 28'b1111111111111110101110101100, 28'b0000000000000000000000000000, 28'b1111111111111111010011110011, 28'b0000000000000000001110101011, 28'b1111111111111100101110110011, 28'b1111111111111111111111111111, 28'b1111111111111111111111110001, 28'b0000000000000001000110011100, 28'b0000000000000010010000001000, 28'b1111111111111101001110000111, 28'b0000000000000010000101001011, 28'b0000000000000000001001011111, 28'b1111111111111111101100111010}, 
{28'b0000000000000001001001101011, 28'b0000000000000100111101100001, 28'b0000000000000001111110110110, 28'b0000000000000001001001000000, 28'b1111111111111110000101101110, 28'b1111111111111110101110101110, 28'b1111111111110101100110100010, 28'b1111111111111110001011000001, 28'b0000000000000001100111001010, 28'b1111111111111111111111111110, 28'b0000000000000001001011010010, 28'b0000000000000011011100111111, 28'b0000000000000000010001110011, 28'b0000000000000000000001011010, 28'b1111111111111111111011101010, 28'b0000000000000000000000000010, 28'b1111111111111111001111100000, 28'b1111111111111111001100001001, 28'b0000000000000000111010111010, 28'b1111111111111101111111011111, 28'b1111111111111101010101110001, 28'b1111111111111111100101101110, 28'b1111111111111101101010100000, 28'b0000000000000000000111100010, 28'b1111111111110110111001001101, 28'b0000000000000011010000101111, 28'b0000000000000011111101001110, 28'b0000000000000010011010100001, 28'b1111111111111001000001101100, 28'b1111111111111110101111111011, 28'b1111111111111101001111111000, 28'b1111111111111100101000000010, 28'b1111111111110101111001100100, 28'b0000000000000010101101001011, 28'b1111111111111111110100110011, 28'b0000000000000001010001100111, 28'b0000000000000000000110000100, 28'b1111111111111010010001001010, 28'b0000000000000000000000000100, 28'b0000000000000000000000000001, 28'b0000000000000000001000001010, 28'b0000000000000100000100111100, 28'b1111111111111111001011100001, 28'b1111111111111101011010111010, 28'b0000000000000011100101101111, 28'b1111111111111110001110011001, 28'b1111111111111110101100111101, 28'b1111111111111110011011100001, 28'b0000000000000001111010001110, 28'b0000000000000010001000000000, 28'b1111111111111111101110100110, 28'b1111111111111110100110101001, 28'b1111111111111111111111011101, 28'b1111111111111111100011001111, 28'b0000000000000000000000000001, 28'b1111111111111110011111011100, 28'b0000000000000010011011010001, 28'b0000000000000100010101100100, 28'b0000000000000010110110001010, 28'b1111111111111100010111010100, 28'b1111111111110001001100000000, 28'b0000000000000011100010101010, 28'b0000000000000000010111101010, 28'b0000000000000001010001001000}, 
{28'b1111111111111111000010001010, 28'b0000000000000001010110010110, 28'b0000000000000001010001010011, 28'b1111111111111111111111100110, 28'b1111111111111110100000110010, 28'b1111111111111111101001000010, 28'b1111111111111110011101110010, 28'b1111111111111111110001110000, 28'b0000000000000000100110001010, 28'b1111111111111111101100110010, 28'b1111111111111111111000000101, 28'b1111111111111111110101111110, 28'b1111111111111111111111110100, 28'b1111111111111111010001000100, 28'b1111111111111111111001001011, 28'b1111111111111111100110010100, 28'b0000000000000001010000001111, 28'b1111111111111111111111111111, 28'b1111111111111101011011111001, 28'b0000000000000001110111000011, 28'b0000000000000010011000011011, 28'b0000000000000001101010001001, 28'b1111111111111110101110110101, 28'b1111111111111111011100111011, 28'b1111111111111110100111011100, 28'b1111111111111110110101110011, 28'b0000000000000000111010000111, 28'b0000000000000000111011111000, 28'b0000000000000000111001111000, 28'b0000000000000001011100000111, 28'b0000000000000000001000110000, 28'b0000000000000001100010110101, 28'b1111111111111111110101010010, 28'b0000000000000000000001001111, 28'b0000000000000001001101111111, 28'b0000000000000000100001101011, 28'b1111111111111111101111000110, 28'b1111111111111111111101100100, 28'b0000000000000000000000000001, 28'b1111111111111110110101000110, 28'b1111111111111111000110110101, 28'b1111111111111111100011110000, 28'b1111111111111110100100000101, 28'b0000000000000001110011001001, 28'b0000000000000000000000000100, 28'b1111111111111111111110100101, 28'b1111111111111111101010110110, 28'b1111111111111111011010001101, 28'b1111111111111100110001110001, 28'b1111111111111111110110000100, 28'b1111111111111111000110100011, 28'b1111111111111111011011101110, 28'b1111111111111111100110011011, 28'b0000000000000001000011101101, 28'b0000000000000010101110100110, 28'b0000000000000000101111111111, 28'b1111111111111111111100100110, 28'b1111111111111110101000001101, 28'b1111111111111111111000011110, 28'b0000000000000000000000000101, 28'b0000000000000001010011010111, 28'b1111111111111111111010100101, 28'b0000000000000000001011101111, 28'b0000000000000000000000000000}
};

localparam logic signed [27:0] bias [64] = '{
28'b1111111111111111110110011100,  // -0.037350185215473175
28'b0000000000000001000110000001,  // 0.27355897426605225
28'b1111111111111111100000010011,  // -0.12378914654254913
28'b1111111111111111101111011111,  // -0.064457006752491
28'b0000000000000000001101111101,  // 0.05452875792980194
28'b0000000000000000011101111000,  // 0.11671770364046097
28'b0000000000000000100010111010,  // 0.13640816509723663
28'b0000000000000000010011001001,  // 0.07482525706291199
28'b0000000000000000001011111101,  // 0.04674031585454941
28'b1111111111111111001100011011,  // -0.20146161317825317
28'b1111111111111111100110101000,  // -0.09910125285387039
28'b0000000000000000100110101010,  // 0.15104414522647858
28'b1111111111111111100101110101,  // -0.10221704095602036
28'b1111111111111111011010100101,  // -0.1461549550294876
28'b1111111111111111101001111000,  // -0.08641516417264938
28'b0000000000000000101010100001,  // 0.16613510251045227
28'b1111111111111111101010100101,  // -0.0836295336484909
28'b1111111111111111110001010000,  // -0.05756539851427078
28'b1111111111111111110111101110,  // -0.03229188174009323
28'b1111111111111111111000101110,  // -0.028388574719429016
28'b0000000000000000100000010000,  // 0.1260243058204651
28'b1111111111111111110110100000,  // -0.037064336240291595
28'b0000000000000000110001100000,  // 0.19336333870887756
28'b0000000000000000000101011100,  // 0.02124214917421341
28'b0000000000000001111111101000,  // 0.4985624849796295
28'b0000000000000000000100000011,  // 0.0158411655575037
28'b1111111111111111101010110000,  // -0.08296407759189606
28'b0000000000000000011100010011,  // 0.11056788265705109
28'b0000000000000000000011000000,  // 0.01173810102045536
28'b1111111111111111100100001111,  // -0.10843746364116669
28'b0000000000000001000110001111,  // 0.27439257502555847
28'b0000000000000000010111100011,  // 0.09199801832437515
28'b0000000000000001000110001100,  // 0.27419957518577576
28'b0000000000000001000101010010,  // 0.27063727378845215
28'b1111111111111111000000011100,  // -0.24828937649726868
28'b0000000000000000010100000000,  // 0.07818280160427094
28'b1111111111111111111110100001,  // -0.005749030504375696
28'b0000000000000000011011110001,  // 0.10850494354963303
28'b0000000000000000100010110010,  // 0.13591453433036804
28'b1111111111111111100001000011,  // -0.12088628858327866
28'b1111111111111111110001011111,  // -0.05666546896100044
28'b0000000000000000010111110101,  // 0.09311636537313461
28'b0000000000000000001110000001,  // 0.05477767437696457
28'b0000000000000000000111100100,  // 0.029585206881165504
28'b1111111111111110110000000110,  // -0.31209176778793335
28'b1111111111111111101010010101,  // -0.08465463668107986
28'b1111111111111111010101000011,  // -0.16775836050510406
28'b0000000000000000100101110010,  // 0.14762157201766968
28'b1111111111111111000011100010,  // -0.23618532717227936
28'b0000000000000000010000101110,  // 0.06535740196704865
28'b1111111111111111011111000110,  // -0.12853026390075684
28'b1111111111111111011100101010,  // -0.13802281022071838
28'b1111111111111111011001001100,  // -0.15156887471675873
28'b0000000000000000010100011011,  // 0.07979883998632431
28'b0000000000000000101110011100,  // 0.18141601979732513
28'b1111111111111111110010001010,  // -0.054039113223552704
28'b1111111111111111111101011011,  // -0.010052933357656002
28'b0000000000000000010000111011,  // 0.06611225008964539
28'b0000000000000000001100111011,  // 0.05053366720676422
28'b0000000000000000000110111000,  // 0.026860840618610382
28'b0000000000000000001000011001,  // 0.03283466026186943
28'b0000000000000000100111110101,  // 0.15558314323425293
28'b1111111111111110110110101100,  // -0.2863388657569885
28'b1111111111111111101001100011   // -0.08769102394580841
};
endpackage