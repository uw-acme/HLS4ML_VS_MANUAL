// Width: 15
// NFRAC: 7
package dense_3_15_7;

localparam logic signed [14:0] weights [32][32] = '{ 
{15'b111111111111001, 15'b111111111001000, 15'b111111111001100, 15'b111111111100111, 15'b000000000101011, 15'b000000000000101, 15'b111111111111110, 15'b111111111111111, 15'b111111111111111, 15'b111111111111111, 15'b000000000010000, 15'b111111110111100, 15'b111111111111000, 15'b000000001101100, 15'b111111111100001, 15'b111111110001000, 15'b111111111111011, 15'b000000000001110, 15'b000000000110111, 15'b111111111010011, 15'b111111101110111, 15'b111111111111010, 15'b000000000000110, 15'b111111111001100, 15'b000000000000000, 15'b000000010000001, 15'b111111101000101, 15'b111111111100011, 15'b111111111001110, 15'b111111111101100, 15'b000000000110110, 15'b111111111101011}, 
{15'b000000001011111, 15'b000000011011101, 15'b000000000110011, 15'b111111110101011, 15'b000000000011111, 15'b111111111011101, 15'b111111111110010, 15'b000000010001011, 15'b000000000000000, 15'b111111111111111, 15'b111111111111011, 15'b111111110110100, 15'b111111111100110, 15'b000000001000101, 15'b111111011110010, 15'b111111111000011, 15'b111111111111111, 15'b111111111111110, 15'b111111111111001, 15'b111111111101010, 15'b111111111011110, 15'b111111111011100, 15'b000000000000010, 15'b111111111111111, 15'b111111111111111, 15'b111111101110110, 15'b000000000000001, 15'b000000000111100, 15'b111111111110111, 15'b111111110100111, 15'b000000000000000, 15'b000000000000100}, 
{15'b111111110000001, 15'b000000000010111, 15'b000000000000001, 15'b000000000101001, 15'b111111110101111, 15'b000000000000000, 15'b000000000000000, 15'b111111110010100, 15'b000000001000100, 15'b111111111011110, 15'b111111111011110, 15'b111111101000001, 15'b111111111011000, 15'b000000001000001, 15'b000000000100001, 15'b111111111111111, 15'b111111111110001, 15'b111111111111100, 15'b111111110010111, 15'b000000000000000, 15'b000000000001111, 15'b000000000001000, 15'b000000000011010, 15'b000000001110000, 15'b000000000000100, 15'b111111110011011, 15'b000000001100010, 15'b000000000000000, 15'b000000000010101, 15'b111111111111101, 15'b000000000000000, 15'b000000100100010}, 
{15'b000000001101011, 15'b111111111111111, 15'b111111111100111, 15'b000000010100111, 15'b000000010011101, 15'b000000000000000, 15'b000000000001001, 15'b000000001101000, 15'b111111111001101, 15'b111111111111111, 15'b111111110010110, 15'b000000000001111, 15'b000000000100010, 15'b111111110100000, 15'b000000000001011, 15'b111111111101011, 15'b111111111111111, 15'b111111111010001, 15'b000000000000100, 15'b000000000000111, 15'b000000000000010, 15'b111111111110110, 15'b000000010011000, 15'b000000001010111, 15'b000000001010100, 15'b000000000111111, 15'b000000001010111, 15'b000000000000000, 15'b111111111110000, 15'b000000001110011, 15'b000000000111111, 15'b111111111101001}, 
{15'b000000010000000, 15'b111111111110100, 15'b111111110100111, 15'b111111100111111, 15'b000000001111010, 15'b000000000000000, 15'b111111110010110, 15'b111111110110111, 15'b111111111110100, 15'b111111100110000, 15'b111111011100101, 15'b000000001111001, 15'b000000010101011, 15'b000000010000101, 15'b111111101101100, 15'b111111100111001, 15'b000000000000000, 15'b111111111011011, 15'b000000000110011, 15'b000000000100011, 15'b111111111001111, 15'b111111111111110, 15'b000000010111000, 15'b111111010100000, 15'b000000000010110, 15'b111111101010111, 15'b000000000010000, 15'b111111111000000, 15'b111111110110011, 15'b111111111111111, 15'b000000000010001, 15'b000000010010100}, 
{15'b000000000001011, 15'b111111111110101, 15'b111111110110001, 15'b111111110111101, 15'b000000001011111, 15'b000000000000000, 15'b111111110111000, 15'b111111111011101, 15'b111111110010010, 15'b111111111101111, 15'b111111111111111, 15'b000000000101001, 15'b000000000000000, 15'b000000001011011, 15'b111111101111110, 15'b111111111011111, 15'b000000000010110, 15'b111111110110100, 15'b111111111001101, 15'b111111111111111, 15'b000000000000011, 15'b000000001001100, 15'b000000001110111, 15'b111111111111101, 15'b111111111111111, 15'b000000001100110, 15'b111111101110011, 15'b111111111111111, 15'b111111111000011, 15'b111111111110110, 15'b111111111111111, 15'b000000000000001}, 
{15'b000000000010000, 15'b111111110101010, 15'b000000000011011, 15'b111111111110110, 15'b111111111111110, 15'b000000000100110, 15'b111111111100100, 15'b111111101010010, 15'b111111111111111, 15'b111111111001010, 15'b111111110001011, 15'b000000001111000, 15'b000000000000001, 15'b000000010101111, 15'b000000011010100, 15'b000000000000000, 15'b111111111111111, 15'b111111110101111, 15'b111111111110000, 15'b000000001000101, 15'b111111100111111, 15'b000000000100111, 15'b000000001010011, 15'b000000000000100, 15'b000000000100110, 15'b000000100111110, 15'b111111110011011, 15'b111111111101000, 15'b111111111001111, 15'b000000001111100, 15'b111111111110011, 15'b111111111010100}, 
{15'b111111101100111, 15'b000000000000110, 15'b111111101011110, 15'b000000001101111, 15'b000000100000111, 15'b000000000011101, 15'b000000000000000, 15'b000000000001100, 15'b111111111111111, 15'b000000000100000, 15'b000000101001101, 15'b111111111111111, 15'b000000001100001, 15'b000000010011111, 15'b000000011000100, 15'b000000100001100, 15'b000000000000000, 15'b111111110000101, 15'b000000001010110, 15'b111111111111110, 15'b111111101011100, 15'b111111111000101, 15'b000000000000011, 15'b111111111101010, 15'b111111101111111, 15'b000000111100000, 15'b111111111000111, 15'b000000000000000, 15'b000000000000000, 15'b000000011100010, 15'b000000000010110, 15'b000000001100100}, 
{15'b000000001101100, 15'b111111111111011, 15'b000000000000000, 15'b111111111110100, 15'b000000000010100, 15'b111111111110110, 15'b111111111111111, 15'b000000000101000, 15'b000000000110110, 15'b111111110111001, 15'b000000000100011, 15'b000000000101111, 15'b000000000000011, 15'b000000001010101, 15'b111111111000110, 15'b111111100110011, 15'b000000000000000, 15'b111111111111100, 15'b111111111111001, 15'b111111110000000, 15'b111111111111111, 15'b000000000000000, 15'b111111111001100, 15'b111111111111100, 15'b111111111100111, 15'b000000000100111, 15'b000000001011111, 15'b111111111100001, 15'b111111111110011, 15'b111111111110101, 15'b000000000000110, 15'b111111110011011}, 
{15'b111111111010010, 15'b000000001100010, 15'b000000000000000, 15'b000000000000000, 15'b000000011001010, 15'b000000001010010, 15'b111111111111111, 15'b111111101110001, 15'b000000000011110, 15'b111111101001101, 15'b111111010011000, 15'b111111111111111, 15'b000000000000000, 15'b000000001101101, 15'b000000000011100, 15'b000000000000000, 15'b111111110101011, 15'b000000000000000, 15'b000000000000001, 15'b000000000001111, 15'b000000000111110, 15'b111111111111001, 15'b111111110100011, 15'b000000000000010, 15'b111111111111101, 15'b000000100010100, 15'b000000001010011, 15'b111111111111111, 15'b111111111101101, 15'b000000010101011, 15'b111111111110101, 15'b111111111101001}, 
{15'b111111101111010, 15'b000000000101100, 15'b111111111110111, 15'b111111111111111, 15'b111111111000000, 15'b111111110011111, 15'b000000000001100, 15'b000000000100100, 15'b111111111111111, 15'b111111111010100, 15'b111111101101101, 15'b000000000110011, 15'b000000001001101, 15'b000000000000000, 15'b000000011010110, 15'b111111101110000, 15'b000000000011010, 15'b111111110011011, 15'b000000001001000, 15'b111111111111111, 15'b111111111110110, 15'b000000000010001, 15'b000000000011111, 15'b000000000000000, 15'b111111110000001, 15'b000000000000111, 15'b111111101110000, 15'b111111111110101, 15'b111111111111111, 15'b000000010101100, 15'b111111111001111, 15'b000000000000000}, 
{15'b111111111111111, 15'b000000000011101, 15'b000000000000000, 15'b000000001100100, 15'b111111111100010, 15'b111111111110100, 15'b000000000001110, 15'b111111111111110, 15'b111111111110100, 15'b000000010100100, 15'b000000010110010, 15'b000000000000000, 15'b111111110101010, 15'b111111101001100, 15'b111111111110011, 15'b000000000000000, 15'b000000000000000, 15'b111111111101111, 15'b111111110000110, 15'b000000001100001, 15'b000000000000000, 15'b000000001011110, 15'b111111111111111, 15'b000000010001111, 15'b000000000011111, 15'b000000001001110, 15'b000000001110100, 15'b111111111110010, 15'b111111110011011, 15'b111111110001111, 15'b111111111111110, 15'b111111101010100}, 
{15'b111111111000110, 15'b111111111111111, 15'b000000000011110, 15'b111111110010100, 15'b000000000010110, 15'b111111111111111, 15'b111111111001000, 15'b111111111111101, 15'b111111111011111, 15'b000000000001001, 15'b000000000010011, 15'b111111111101101, 15'b000000000000100, 15'b000000000110000, 15'b111111101011111, 15'b111111111000001, 15'b000000000111010, 15'b111111111010010, 15'b000000000000000, 15'b111111111111001, 15'b000000000110001, 15'b000000000000010, 15'b111111111111000, 15'b000000000001010, 15'b000000001000100, 15'b111111111100101, 15'b000000000000000, 15'b111111110001100, 15'b111111111001101, 15'b111111111111110, 15'b000000000101100, 15'b000000000000000}, 
{15'b111111101111010, 15'b000000001101011, 15'b111111111111111, 15'b111111111111110, 15'b111111111111101, 15'b000000000101100, 15'b111111111111111, 15'b000000011000101, 15'b111111111111100, 15'b111111111111111, 15'b000000000110100, 15'b000000000001010, 15'b000000000000001, 15'b000000000000000, 15'b000000000011111, 15'b000000001010100, 15'b000000000101101, 15'b000000000101010, 15'b111111111111101, 15'b000000001001110, 15'b000000000011001, 15'b000000000001010, 15'b111111111111101, 15'b000000001000001, 15'b111111111100110, 15'b111111110101001, 15'b111111111101000, 15'b111111111111111, 15'b000000000011010, 15'b000000000000111, 15'b000000000110010, 15'b000000001111010}, 
{15'b111111111111011, 15'b111111110011100, 15'b000000000001101, 15'b111111111111111, 15'b000000011101010, 15'b111111111001010, 15'b111111101101101, 15'b000000000000000, 15'b000000000000000, 15'b111111111111001, 15'b000000000001100, 15'b000000001101111, 15'b000000001010010, 15'b000000000000010, 15'b000000000001000, 15'b111111111010011, 15'b000000000001000, 15'b111111111110110, 15'b000000000000000, 15'b000000000010011, 15'b111111111110110, 15'b000000000000100, 15'b000000001000100, 15'b000000000001001, 15'b111111111111100, 15'b111111110010110, 15'b000000000110100, 15'b111111111111111, 15'b111111111111111, 15'b111111111100100, 15'b111111111111010, 15'b111111111101111}, 
{15'b000000000000001, 15'b111111111101111, 15'b111111111011111, 15'b111111111001000, 15'b111111101110100, 15'b000000010011100, 15'b000000000000000, 15'b000000000101011, 15'b000000001001001, 15'b000000000000011, 15'b111111111110111, 15'b000000001111001, 15'b000000000111001, 15'b111111110100010, 15'b111111111010110, 15'b111111111110101, 15'b111111110011010, 15'b111111111111011, 15'b000000000000000, 15'b111111111111110, 15'b000000000100111, 15'b111111111011100, 15'b000000000000000, 15'b000000000010011, 15'b111111111111111, 15'b111111110101000, 15'b000000000101000, 15'b000000000000000, 15'b000000000001011, 15'b000000000000010, 15'b111111110101111, 15'b000000000000101}, 
{15'b111111111001101, 15'b111111111010111, 15'b000000000010011, 15'b111111111100000, 15'b111111111101001, 15'b000000000011101, 15'b111111111111110, 15'b000000000001000, 15'b000000000100001, 15'b111111111111111, 15'b000000000011111, 15'b111111111011111, 15'b111111111111101, 15'b111111111111111, 15'b000000000011010, 15'b111111111111111, 15'b000000001111101, 15'b111111111111011, 15'b000000000111111, 15'b111111111010100, 15'b000000000101000, 15'b000000000010000, 15'b000000000010101, 15'b000000000001001, 15'b111111111101011, 15'b111111110111000, 15'b111111110111101, 15'b000000000011011, 15'b111111111101010, 15'b000000000000000, 15'b111111111111000, 15'b000000000111011}, 
{15'b111111111111111, 15'b111111110011000, 15'b111111110011010, 15'b111111111111111, 15'b000000010100001, 15'b111111111101000, 15'b000000000000000, 15'b000000001111011, 15'b111111111011010, 15'b000000000000000, 15'b111111110010101, 15'b111111110000010, 15'b000000001110010, 15'b000000000100110, 15'b111111111100000, 15'b111111110111001, 15'b000000000101100, 15'b000000000000000, 15'b111111111000011, 15'b000000000000110, 15'b000000000010001, 15'b111111111101001, 15'b000000001001000, 15'b111111100000101, 15'b000000000001010, 15'b000000000111101, 15'b111111111110101, 15'b000000000000011, 15'b111111111000100, 15'b111111111111111, 15'b111111111001100, 15'b111111111111001}, 
{15'b000000000110110, 15'b000000001011000, 15'b000000010001100, 15'b111111111001011, 15'b000000001101010, 15'b000000001001110, 15'b000000000000000, 15'b000000001110100, 15'b000000001011011, 15'b111111111100100, 15'b000000010110011, 15'b111111110100110, 15'b000000010011111, 15'b000000001110010, 15'b111111011101101, 15'b111111111111111, 15'b000000000000000, 15'b000000000000001, 15'b000000001000010, 15'b111111101111111, 15'b000000000111000, 15'b111111111001001, 15'b111111110000010, 15'b111111111010111, 15'b000000001010100, 15'b111111101010111, 15'b111111110101011, 15'b111111111110101, 15'b111111111111111, 15'b111111101101111, 15'b000000001100101, 15'b000000000000000}, 
{15'b111111111110011, 15'b000000000000000, 15'b111111111111111, 15'b111111111111111, 15'b111111110100110, 15'b000000000000010, 15'b000000000000010, 15'b111111111111100, 15'b111111111111001, 15'b111111111110100, 15'b000000000100011, 15'b111111111111111, 15'b000000000010101, 15'b111111110101000, 15'b000000000011011, 15'b111111111111111, 15'b000000000100100, 15'b000000001110010, 15'b111111110100101, 15'b000000000001101, 15'b111111111100110, 15'b000000000100000, 15'b000000000110000, 15'b111111111101010, 15'b111111110111111, 15'b000000000000101, 15'b000000011010100, 15'b111111111111001, 15'b111111111111100, 15'b000000001010011, 15'b000000000000000, 15'b000000011011100}, 
{15'b111111101111010, 15'b000000000001001, 15'b111111111001000, 15'b000000001100010, 15'b000000000011100, 15'b111111111110111, 15'b111111111111111, 15'b111111111111111, 15'b111111110110010, 15'b111111111110111, 15'b000000000000000, 15'b111111101110001, 15'b000000000000011, 15'b111111111110101, 15'b111111111111111, 15'b111111111111111, 15'b111111111100010, 15'b000000000000001, 15'b000000000000000, 15'b000000000101000, 15'b000000000000100, 15'b000000000000000, 15'b000000000000000, 15'b111111111111101, 15'b000000000000000, 15'b000000000000100, 15'b000000010010100, 15'b111111111111111, 15'b111111111111111, 15'b111111111110101, 15'b000000000101100, 15'b111111111111001}, 
{15'b111111111111111, 15'b111111111011001, 15'b000000000110100, 15'b000000000001010, 15'b111111110100000, 15'b000000000000000, 15'b000000001001001, 15'b111111111111111, 15'b000000000000000, 15'b111111111100110, 15'b000000000011101, 15'b000000000000100, 15'b000000001010010, 15'b111111101110011, 15'b111111111100111, 15'b111111111111011, 15'b000000000110111, 15'b111111110011101, 15'b000000000000101, 15'b111111100111110, 15'b111111111111011, 15'b111111111100001, 15'b111111111110101, 15'b000000001001011, 15'b111111111101100, 15'b111111110111000, 15'b000000000010111, 15'b000000000000000, 15'b000000001100101, 15'b000000010000101, 15'b111111110101100, 15'b111111110001101}, 
{15'b000000000010001, 15'b000000000000110, 15'b111111110010101, 15'b111111111110001, 15'b111111111111111, 15'b000000000000000, 15'b000000000011011, 15'b000000001101001, 15'b000000000000000, 15'b000000000000101, 15'b000000000010001, 15'b111111101110101, 15'b111111111101110, 15'b111111101100101, 15'b000000001111011, 15'b000000000000000, 15'b111111111111111, 15'b111111101011011, 15'b111111111111111, 15'b111111111101100, 15'b111111111111010, 15'b000000000000000, 15'b000000000001111, 15'b111111111011001, 15'b000000000001101, 15'b000000001101001, 15'b000000001101101, 15'b000000001100011, 15'b000000001001110, 15'b000000000000000, 15'b000000000011101, 15'b000000011001000}, 
{15'b111111111111001, 15'b111111111000011, 15'b000000001100011, 15'b111111111100101, 15'b000000000010001, 15'b000000000101010, 15'b111111111111111, 15'b111111110110110, 15'b111111111101010, 15'b111111101100110, 15'b000000001110010, 15'b000000000000000, 15'b000000001101011, 15'b000000010101011, 15'b111111111100010, 15'b111111100100001, 15'b111111111100101, 15'b000000001111000, 15'b111111110110111, 15'b111111111001010, 15'b000000000001111, 15'b000000000000000, 15'b111111101110100, 15'b111111111001111, 15'b111111111110101, 15'b111111111100000, 15'b000000000011100, 15'b000000010110100, 15'b000000000111110, 15'b111111111111111, 15'b000000000010100, 15'b000000000000111}, 
{15'b000000000001010, 15'b000000001110100, 15'b000000000000000, 15'b000000001001011, 15'b000000011010100, 15'b111111111010100, 15'b111111111111111, 15'b111111111110100, 15'b000000001001011, 15'b111111111001110, 15'b111111111111111, 15'b000000001010101, 15'b000000000000010, 15'b000000000000111, 15'b111111001111001, 15'b111111111101011, 15'b000000000000000, 15'b000000000110011, 15'b111111111111111, 15'b000000001001100, 15'b111111111111111, 15'b111111111010011, 15'b111111101110000, 15'b000000000100001, 15'b000000001001001, 15'b111111011100100, 15'b111111111111111, 15'b000000000000000, 15'b000000010001011, 15'b111111100110010, 15'b000000000000000, 15'b111111111111110}, 
{15'b000000000000010, 15'b111111110101001, 15'b000000000001101, 15'b111111111111100, 15'b000000000001101, 15'b000000010000111, 15'b111111101000110, 15'b000000000001000, 15'b000000001101100, 15'b111111110101001, 15'b111111111111010, 15'b000000000001100, 15'b111111111111101, 15'b000000000101101, 15'b000000000011011, 15'b111111111111011, 15'b000000000010001, 15'b000000000000000, 15'b000000000000101, 15'b000000001100001, 15'b111111111111000, 15'b111111110000100, 15'b111111101100101, 15'b111111111001110, 15'b111111101101000, 15'b000000000110101, 15'b000000010011111, 15'b000000001011110, 15'b111111111111101, 15'b111111110100000, 15'b111111110110000, 15'b000000000001111}, 
{15'b000000000001101, 15'b111111110000101, 15'b111111111111011, 15'b000000000100110, 15'b111111110000101, 15'b000000000101011, 15'b111111111111111, 15'b111111111111111, 15'b111111111111111, 15'b000000000000000, 15'b000000001000011, 15'b111111111111011, 15'b000000000000010, 15'b000000000000000, 15'b000000000100000, 15'b111111111111011, 15'b000000000000000, 15'b111111111111111, 15'b111111110101101, 15'b111111101111110, 15'b111111111111111, 15'b111111101110111, 15'b111111110110010, 15'b111111110100000, 15'b000000011100011, 15'b000000000000100, 15'b111111111110100, 15'b000000001010001, 15'b000000011100101, 15'b000000001100101, 15'b111111011110000, 15'b111111111010000}, 
{15'b000000001100000, 15'b111111111111111, 15'b000000001000000, 15'b111111111111010, 15'b000000001111011, 15'b111111111011011, 15'b000000000010010, 15'b000000001101011, 15'b000000001000100, 15'b111111101111010, 15'b111111111110000, 15'b000000000011111, 15'b000000000010001, 15'b111111111111100, 15'b000000000010101, 15'b000000000000000, 15'b000000001011100, 15'b000000000001000, 15'b000000001011111, 15'b111111111101111, 15'b111111111011111, 15'b111111111101100, 15'b111111111111111, 15'b000000001001101, 15'b111111111001100, 15'b111111111111110, 15'b000000000000000, 15'b000000000000000, 15'b000000000000000, 15'b000000001001010, 15'b111111110101101, 15'b111111111111010}, 
{15'b111111111111111, 15'b111111111111000, 15'b111111110001000, 15'b000000001001000, 15'b000000000111001, 15'b111111111100011, 15'b111111111111111, 15'b111111111000101, 15'b000000000000001, 15'b111111111111111, 15'b111111110110010, 15'b111111111000000, 15'b000000001111010, 15'b000000000000000, 15'b111111111011111, 15'b111111111111111, 15'b000000000110110, 15'b111111111111111, 15'b111111111111111, 15'b111111111001000, 15'b000000001010000, 15'b000000000000000, 15'b000000000100111, 15'b111111111111000, 15'b000000000101000, 15'b000000000000000, 15'b000000000000000, 15'b000000000111101, 15'b111111111001110, 15'b111111111110100, 15'b000000000101001, 15'b111111111100100}, 
{15'b111111111111011, 15'b111111110110001, 15'b000000010011000, 15'b111111111101111, 15'b000000000110010, 15'b111111110110110, 15'b000000000000000, 15'b000000000001000, 15'b111111110000101, 15'b111111111111100, 15'b111111111100000, 15'b000000000001110, 15'b111111110101100, 15'b000000000100011, 15'b000000000110011, 15'b000000000011100, 15'b000000000010101, 15'b111111111110110, 15'b111111101001010, 15'b111111111111100, 15'b111111111110001, 15'b000000000100011, 15'b111111111100011, 15'b111111111111111, 15'b000000000110010, 15'b111111111110100, 15'b111111111111100, 15'b000000001100011, 15'b111111110011010, 15'b111111110110100, 15'b000000001011001, 15'b000000000001001}, 
{15'b000000001101110, 15'b000000000110011, 15'b000000000000000, 15'b111111111010111, 15'b111111111101011, 15'b111111111111111, 15'b000000000000000, 15'b111111111101110, 15'b111111111100000, 15'b111111111100001, 15'b000000000000000, 15'b000000000101000, 15'b000000000000001, 15'b000000000001101, 15'b111111111110100, 15'b000000000000001, 15'b111111111011000, 15'b000000000000000, 15'b111111111111011, 15'b111111111111111, 15'b000000000000000, 15'b000000000001111, 15'b000000000011000, 15'b000000000000000, 15'b000000000000000, 15'b111111101100011, 15'b111111111001100, 15'b000000000000001, 15'b000000000000101, 15'b000000000000000, 15'b111111111010010, 15'b000000000000101}, 
{15'b000000000110000, 15'b111111011110100, 15'b111111111111111, 15'b111111111101100, 15'b111111111000100, 15'b111111111111101, 15'b000000000000000, 15'b000000010001100, 15'b111111111110100, 15'b111111111111010, 15'b000000000010101, 15'b111111101010110, 15'b000000000000110, 15'b111111110001111, 15'b000000010111000, 15'b111111111110010, 15'b111111111000110, 15'b111111101110011, 15'b111111111111101, 15'b111111101001010, 15'b111111100110000, 15'b111111111111111, 15'b000000000000000, 15'b000000000000000, 15'b000000000111110, 15'b111111111111100, 15'b111111110110011, 15'b111111111101101, 15'b111111111111010, 15'b000000000000000, 15'b111111111110111, 15'b111111101001100}
};

localparam logic signed [14:0] bias [32] = '{
15'b000000001000011,  // 0.5280959606170654
15'b000000001101011,  // 0.8414360880851746
15'b000000000110010,  // 0.397830605506897
15'b000000000110100,  // 0.4105983078479767
15'b111111000101011,  // -3.657735586166382
15'b111111110001101,  // -0.8977976441383362
15'b000000011011010,  // 1.7051936388015747
15'b111111101011100,  // -1.2765135765075684
15'b111111110110101,  // -0.5837795734405518
15'b000000101011001,  // 2.699671983718872
15'b000000000011011,  // 0.2170683741569519
15'b000000001110000,  // 0.8814588785171509
15'b111111010101110,  // -2.634300947189331
15'b111111100001111,  // -1.877297282218933
15'b000000011010100,  // 1.6625694036483765
15'b000000101011111,  // 2.7459704875946045
15'b111111111000010,  // -0.47838035225868225
15'b000000011011001,  // 1.6984987258911133
15'b000000001101101,  // 0.8548859357833862
15'b000000010000000,  // 1.0045719146728516
15'b000000010110101,  // 1.4197649955749512
15'b000000001101010,  // 0.832463800907135
15'b000000001000101,  // 0.5434179306030273
15'b000000001110110,  // 0.9277304410934448
15'b111111111010100,  // -0.3426123857498169
15'b111111110111000,  // -0.5587119460105896
15'b111111110110000,  // -0.6208624839782715
15'b111111101011100,  // -1.2802538871765137
15'b000000000000111,  // 0.05940237268805504
15'b111111110010110,  // -0.8213341236114502
15'b000000001110000,  // 0.8783953189849854
15'b111111110000110   // -0.949700653553009
};
endpackage