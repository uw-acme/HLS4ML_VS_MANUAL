// Width: 10
// NFRAC: 5
package dense_3_10_5;

localparam logic signed [9:0] weights [32][32] = '{ 
{10'b1111111110, 10'b1111110010, 10'b1111110011, 10'b1111111001, 10'b0000001010, 10'b0000000001, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b0000000100, 10'b1111101111, 10'b1111111110, 10'b0000011011, 10'b1111111000, 10'b1111100010, 10'b1111111110, 10'b0000000011, 10'b0000001101, 10'b1111110100, 10'b1111011101, 10'b1111111110, 10'b0000000001, 10'b1111110011, 10'b0000000000, 10'b0000100000, 10'b1111010001, 10'b1111111000, 10'b1111110011, 10'b1111111011, 10'b0000001101, 10'b1111111010}, 
{10'b0000010111, 10'b0000110111, 10'b0000001100, 10'b1111101010, 10'b0000000111, 10'b1111110111, 10'b1111111100, 10'b0000100010, 10'b0000000000, 10'b1111111111, 10'b1111111110, 10'b1111101101, 10'b1111111001, 10'b0000010001, 10'b1110111100, 10'b1111110000, 10'b1111111111, 10'b1111111111, 10'b1111111110, 10'b1111111010, 10'b1111110111, 10'b1111110111, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b1111011101, 10'b0000000000, 10'b0000001111, 10'b1111111101, 10'b1111101001, 10'b0000000000, 10'b0000000001}, 
{10'b1111100000, 10'b0000000101, 10'b0000000000, 10'b0000001010, 10'b1111101011, 10'b0000000000, 10'b0000000000, 10'b1111100101, 10'b0000010001, 10'b1111110111, 10'b1111110111, 10'b1111010000, 10'b1111110110, 10'b0000010000, 10'b0000001000, 10'b1111111111, 10'b1111111100, 10'b1111111111, 10'b1111100101, 10'b0000000000, 10'b0000000011, 10'b0000000010, 10'b0000000110, 10'b0000011100, 10'b0000000001, 10'b1111100110, 10'b0000011000, 10'b0000000000, 10'b0000000101, 10'b1111111111, 10'b0000000000, 10'b0001001000}, 
{10'b0000011010, 10'b1111111111, 10'b1111111001, 10'b0000101001, 10'b0000100111, 10'b0000000000, 10'b0000000010, 10'b0000011010, 10'b1111110011, 10'b1111111111, 10'b1111100101, 10'b0000000011, 10'b0000001000, 10'b1111101000, 10'b0000000010, 10'b1111111010, 10'b1111111111, 10'b1111110100, 10'b0000000001, 10'b0000000001, 10'b0000000000, 10'b1111111101, 10'b0000100110, 10'b0000010101, 10'b0000010101, 10'b0000001111, 10'b0000010101, 10'b0000000000, 10'b1111111100, 10'b0000011100, 10'b0000001111, 10'b1111111010}, 
{10'b0000100000, 10'b1111111101, 10'b1111101001, 10'b1111001111, 10'b0000011110, 10'b0000000000, 10'b1111100101, 10'b1111101101, 10'b1111111101, 10'b1111001100, 10'b1110111001, 10'b0000011110, 10'b0000101010, 10'b0000100001, 10'b1111011011, 10'b1111001110, 10'b0000000000, 10'b1111110110, 10'b0000001100, 10'b0000001000, 10'b1111110011, 10'b1111111111, 10'b0000101110, 10'b1110101000, 10'b0000000101, 10'b1111010101, 10'b0000000100, 10'b1111110000, 10'b1111101100, 10'b1111111111, 10'b0000000100, 10'b0000100101}, 
{10'b0000000010, 10'b1111111101, 10'b1111101100, 10'b1111101111, 10'b0000010111, 10'b0000000000, 10'b1111101110, 10'b1111110111, 10'b1111100100, 10'b1111111011, 10'b1111111111, 10'b0000001010, 10'b0000000000, 10'b0000010110, 10'b1111011111, 10'b1111110111, 10'b0000000101, 10'b1111101101, 10'b1111110011, 10'b1111111111, 10'b0000000000, 10'b0000010011, 10'b0000011101, 10'b1111111111, 10'b1111111111, 10'b0000011001, 10'b1111011100, 10'b1111111111, 10'b1111110000, 10'b1111111101, 10'b1111111111, 10'b0000000000}, 
{10'b0000000100, 10'b1111101010, 10'b0000000110, 10'b1111111101, 10'b1111111111, 10'b0000001001, 10'b1111111001, 10'b1111010100, 10'b1111111111, 10'b1111110010, 10'b1111100010, 10'b0000011110, 10'b0000000000, 10'b0000101011, 10'b0000110101, 10'b0000000000, 10'b1111111111, 10'b1111101011, 10'b1111111100, 10'b0000010001, 10'b1111001111, 10'b0000001001, 10'b0000010100, 10'b0000000001, 10'b0000001001, 10'b0001001111, 10'b1111100110, 10'b1111111010, 10'b1111110011, 10'b0000011111, 10'b1111111100, 10'b1111110101}, 
{10'b1111011001, 10'b0000000001, 10'b1111010111, 10'b0000011011, 10'b0001000001, 10'b0000000111, 10'b0000000000, 10'b0000000011, 10'b1111111111, 10'b0000001000, 10'b0001010011, 10'b1111111111, 10'b0000011000, 10'b0000100111, 10'b0000110001, 10'b0001000011, 10'b0000000000, 10'b1111100001, 10'b0000010101, 10'b1111111111, 10'b1111010111, 10'b1111110001, 10'b0000000000, 10'b1111111010, 10'b1111011111, 10'b0001111000, 10'b1111110001, 10'b0000000000, 10'b0000000000, 10'b0000111000, 10'b0000000101, 10'b0000011001}, 
{10'b0000011011, 10'b1111111110, 10'b0000000000, 10'b1111111101, 10'b0000000101, 10'b1111111101, 10'b1111111111, 10'b0000001010, 10'b0000001101, 10'b1111101110, 10'b0000001000, 10'b0000001011, 10'b0000000000, 10'b0000010101, 10'b1111110001, 10'b1111001100, 10'b0000000000, 10'b1111111111, 10'b1111111110, 10'b1111100000, 10'b1111111111, 10'b0000000000, 10'b1111110011, 10'b1111111111, 10'b1111111001, 10'b0000001001, 10'b0000010111, 10'b1111111000, 10'b1111111100, 10'b1111111101, 10'b0000000001, 10'b1111100110}, 
{10'b1111110100, 10'b0000011000, 10'b0000000000, 10'b0000000000, 10'b0000110010, 10'b0000010100, 10'b1111111111, 10'b1111011100, 10'b0000000111, 10'b1111010011, 10'b1110100110, 10'b1111111111, 10'b0000000000, 10'b0000011011, 10'b0000000111, 10'b0000000000, 10'b1111101010, 10'b0000000000, 10'b0000000000, 10'b0000000011, 10'b0000001111, 10'b1111111110, 10'b1111101000, 10'b0000000000, 10'b1111111111, 10'b0001000101, 10'b0000010100, 10'b1111111111, 10'b1111111011, 10'b0000101010, 10'b1111111101, 10'b1111111010}, 
{10'b1111011110, 10'b0000001011, 10'b1111111101, 10'b1111111111, 10'b1111110000, 10'b1111100111, 10'b0000000011, 10'b0000001001, 10'b1111111111, 10'b1111110101, 10'b1111011011, 10'b0000001100, 10'b0000010011, 10'b0000000000, 10'b0000110101, 10'b1111011100, 10'b0000000110, 10'b1111100110, 10'b0000010010, 10'b1111111111, 10'b1111111101, 10'b0000000100, 10'b0000000111, 10'b0000000000, 10'b1111100000, 10'b0000000001, 10'b1111011100, 10'b1111111101, 10'b1111111111, 10'b0000101011, 10'b1111110011, 10'b0000000000}, 
{10'b1111111111, 10'b0000000111, 10'b0000000000, 10'b0000011001, 10'b1111111000, 10'b1111111101, 10'b0000000011, 10'b1111111111, 10'b1111111101, 10'b0000101001, 10'b0000101100, 10'b0000000000, 10'b1111101010, 10'b1111010011, 10'b1111111100, 10'b0000000000, 10'b0000000000, 10'b1111111011, 10'b1111100001, 10'b0000011000, 10'b0000000000, 10'b0000010111, 10'b1111111111, 10'b0000100011, 10'b0000000111, 10'b0000010011, 10'b0000011101, 10'b1111111100, 10'b1111100110, 10'b1111100011, 10'b1111111111, 10'b1111010101}, 
{10'b1111110001, 10'b1111111111, 10'b0000000111, 10'b1111100101, 10'b0000000101, 10'b1111111111, 10'b1111110010, 10'b1111111111, 10'b1111110111, 10'b0000000010, 10'b0000000100, 10'b1111111011, 10'b0000000001, 10'b0000001100, 10'b1111010111, 10'b1111110000, 10'b0000001110, 10'b1111110100, 10'b0000000000, 10'b1111111110, 10'b0000001100, 10'b0000000000, 10'b1111111110, 10'b0000000010, 10'b0000010001, 10'b1111111001, 10'b0000000000, 10'b1111100011, 10'b1111110011, 10'b1111111111, 10'b0000001011, 10'b0000000000}, 
{10'b1111011110, 10'b0000011010, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b0000001011, 10'b1111111111, 10'b0000110001, 10'b1111111111, 10'b1111111111, 10'b0000001101, 10'b0000000010, 10'b0000000000, 10'b0000000000, 10'b0000000111, 10'b0000010101, 10'b0000001011, 10'b0000001010, 10'b1111111111, 10'b0000010011, 10'b0000000110, 10'b0000000010, 10'b1111111111, 10'b0000010000, 10'b1111111001, 10'b1111101010, 10'b1111111010, 10'b1111111111, 10'b0000000110, 10'b0000000001, 10'b0000001100, 10'b0000011110}, 
{10'b1111111110, 10'b1111100111, 10'b0000000011, 10'b1111111111, 10'b0000111010, 10'b1111110010, 10'b1111011011, 10'b0000000000, 10'b0000000000, 10'b1111111110, 10'b0000000011, 10'b0000011011, 10'b0000010100, 10'b0000000000, 10'b0000000010, 10'b1111110100, 10'b0000000010, 10'b1111111101, 10'b0000000000, 10'b0000000100, 10'b1111111101, 10'b0000000001, 10'b0000010001, 10'b0000000010, 10'b1111111111, 10'b1111100101, 10'b0000001101, 10'b1111111111, 10'b1111111111, 10'b1111111001, 10'b1111111110, 10'b1111111011}, 
{10'b0000000000, 10'b1111111011, 10'b1111110111, 10'b1111110010, 10'b1111011101, 10'b0000100111, 10'b0000000000, 10'b0000001010, 10'b0000010010, 10'b0000000000, 10'b1111111101, 10'b0000011110, 10'b0000001110, 10'b1111101000, 10'b1111110101, 10'b1111111101, 10'b1111100110, 10'b1111111110, 10'b0000000000, 10'b1111111111, 10'b0000001001, 10'b1111110111, 10'b0000000000, 10'b0000000100, 10'b1111111111, 10'b1111101010, 10'b0000001010, 10'b0000000000, 10'b0000000010, 10'b0000000000, 10'b1111101011, 10'b0000000001}, 
{10'b1111110011, 10'b1111110101, 10'b0000000100, 10'b1111111000, 10'b1111111010, 10'b0000000111, 10'b1111111111, 10'b0000000010, 10'b0000001000, 10'b1111111111, 10'b0000000111, 10'b1111110111, 10'b1111111111, 10'b1111111111, 10'b0000000110, 10'b1111111111, 10'b0000011111, 10'b1111111110, 10'b0000001111, 10'b1111110101, 10'b0000001010, 10'b0000000100, 10'b0000000101, 10'b0000000010, 10'b1111111010, 10'b1111101110, 10'b1111101111, 10'b0000000110, 10'b1111111010, 10'b0000000000, 10'b1111111110, 10'b0000001110}, 
{10'b1111111111, 10'b1111100110, 10'b1111100110, 10'b1111111111, 10'b0000101000, 10'b1111111010, 10'b0000000000, 10'b0000011110, 10'b1111110110, 10'b0000000000, 10'b1111100101, 10'b1111100000, 10'b0000011100, 10'b0000001001, 10'b1111111000, 10'b1111101110, 10'b0000001011, 10'b0000000000, 10'b1111110000, 10'b0000000001, 10'b0000000100, 10'b1111111010, 10'b0000010010, 10'b1111000001, 10'b0000000010, 10'b0000001111, 10'b1111111101, 10'b0000000000, 10'b1111110001, 10'b1111111111, 10'b1111110011, 10'b1111111110}, 
{10'b0000001101, 10'b0000010110, 10'b0000100011, 10'b1111110010, 10'b0000011010, 10'b0000010011, 10'b0000000000, 10'b0000011101, 10'b0000010110, 10'b1111111001, 10'b0000101100, 10'b1111101001, 10'b0000100111, 10'b0000011100, 10'b1110111011, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b0000010000, 10'b1111011111, 10'b0000001110, 10'b1111110010, 10'b1111100000, 10'b1111110101, 10'b0000010101, 10'b1111010101, 10'b1111101010, 10'b1111111101, 10'b1111111111, 10'b1111011011, 10'b0000011001, 10'b0000000000}, 
{10'b1111111100, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b1111101001, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b1111111110, 10'b1111111101, 10'b0000001000, 10'b1111111111, 10'b0000000101, 10'b1111101010, 10'b0000000110, 10'b1111111111, 10'b0000001001, 10'b0000011100, 10'b1111101001, 10'b0000000011, 10'b1111111001, 10'b0000001000, 10'b0000001100, 10'b1111111010, 10'b1111101111, 10'b0000000001, 10'b0000110101, 10'b1111111110, 10'b1111111111, 10'b0000010100, 10'b0000000000, 10'b0000110111}, 
{10'b1111011110, 10'b0000000010, 10'b1111110010, 10'b0000011000, 10'b0000000111, 10'b1111111101, 10'b1111111111, 10'b1111111111, 10'b1111101100, 10'b1111111101, 10'b0000000000, 10'b1111011100, 10'b0000000000, 10'b1111111101, 10'b1111111111, 10'b1111111111, 10'b1111111000, 10'b0000000000, 10'b0000000000, 10'b0000001010, 10'b0000000001, 10'b0000000000, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b0000000001, 10'b0000100101, 10'b1111111111, 10'b1111111111, 10'b1111111101, 10'b0000001011, 10'b1111111110}, 
{10'b1111111111, 10'b1111110110, 10'b0000001101, 10'b0000000010, 10'b1111101000, 10'b0000000000, 10'b0000010010, 10'b1111111111, 10'b0000000000, 10'b1111111001, 10'b0000000111, 10'b0000000001, 10'b0000010100, 10'b1111011100, 10'b1111111001, 10'b1111111110, 10'b0000001101, 10'b1111100111, 10'b0000000001, 10'b1111001111, 10'b1111111110, 10'b1111111000, 10'b1111111101, 10'b0000010010, 10'b1111111011, 10'b1111101110, 10'b0000000101, 10'b0000000000, 10'b0000011001, 10'b0000100001, 10'b1111101011, 10'b1111100011}, 
{10'b0000000100, 10'b0000000001, 10'b1111100101, 10'b1111111100, 10'b1111111111, 10'b0000000000, 10'b0000000110, 10'b0000011010, 10'b0000000000, 10'b0000000001, 10'b0000000100, 10'b1111011101, 10'b1111111011, 10'b1111011001, 10'b0000011110, 10'b0000000000, 10'b1111111111, 10'b1111010110, 10'b1111111111, 10'b1111111011, 10'b1111111110, 10'b0000000000, 10'b0000000011, 10'b1111110110, 10'b0000000011, 10'b0000011010, 10'b0000011011, 10'b0000011000, 10'b0000010011, 10'b0000000000, 10'b0000000111, 10'b0000110010}, 
{10'b1111111110, 10'b1111110000, 10'b0000011000, 10'b1111111001, 10'b0000000100, 10'b0000001010, 10'b1111111111, 10'b1111101101, 10'b1111111010, 10'b1111011001, 10'b0000011100, 10'b0000000000, 10'b0000011010, 10'b0000101010, 10'b1111111000, 10'b1111001000, 10'b1111111001, 10'b0000011110, 10'b1111101101, 10'b1111110010, 10'b0000000011, 10'b0000000000, 10'b1111011101, 10'b1111110011, 10'b1111111101, 10'b1111111000, 10'b0000000111, 10'b0000101101, 10'b0000001111, 10'b1111111111, 10'b0000000101, 10'b0000000001}, 
{10'b0000000010, 10'b0000011101, 10'b0000000000, 10'b0000010010, 10'b0000110101, 10'b1111110101, 10'b1111111111, 10'b1111111101, 10'b0000010010, 10'b1111110011, 10'b1111111111, 10'b0000010101, 10'b0000000000, 10'b0000000001, 10'b1110011110, 10'b1111111010, 10'b0000000000, 10'b0000001100, 10'b1111111111, 10'b0000010011, 10'b1111111111, 10'b1111110100, 10'b1111011100, 10'b0000001000, 10'b0000010010, 10'b1110111001, 10'b1111111111, 10'b0000000000, 10'b0000100010, 10'b1111001100, 10'b0000000000, 10'b1111111111}, 
{10'b0000000000, 10'b1111101010, 10'b0000000011, 10'b1111111111, 10'b0000000011, 10'b0000100001, 10'b1111010001, 10'b0000000010, 10'b0000011011, 10'b1111101010, 10'b1111111110, 10'b0000000011, 10'b1111111111, 10'b0000001011, 10'b0000000110, 10'b1111111110, 10'b0000000100, 10'b0000000000, 10'b0000000001, 10'b0000011000, 10'b1111111110, 10'b1111100001, 10'b1111011001, 10'b1111110011, 10'b1111011010, 10'b0000001101, 10'b0000100111, 10'b0000010111, 10'b1111111111, 10'b1111101000, 10'b1111101100, 10'b0000000011}, 
{10'b0000000011, 10'b1111100001, 10'b1111111110, 10'b0000001001, 10'b1111100001, 10'b0000001010, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b0000000000, 10'b0000010000, 10'b1111111110, 10'b0000000000, 10'b0000000000, 10'b0000001000, 10'b1111111110, 10'b0000000000, 10'b1111111111, 10'b1111101011, 10'b1111011111, 10'b1111111111, 10'b1111011101, 10'b1111101100, 10'b1111101000, 10'b0000111000, 10'b0000000001, 10'b1111111101, 10'b0000010100, 10'b0000111001, 10'b0000011001, 10'b1110111100, 10'b1111110100}, 
{10'b0000011000, 10'b1111111111, 10'b0000010000, 10'b1111111110, 10'b0000011110, 10'b1111110110, 10'b0000000100, 10'b0000011010, 10'b0000010001, 10'b1111011110, 10'b1111111100, 10'b0000000111, 10'b0000000100, 10'b1111111111, 10'b0000000101, 10'b0000000000, 10'b0000010111, 10'b0000000010, 10'b0000010111, 10'b1111111011, 10'b1111110111, 10'b1111111011, 10'b1111111111, 10'b0000010011, 10'b1111110011, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b0000000000, 10'b0000010010, 10'b1111101011, 10'b1111111110}, 
{10'b1111111111, 10'b1111111110, 10'b1111100010, 10'b0000010010, 10'b0000001110, 10'b1111111000, 10'b1111111111, 10'b1111110001, 10'b0000000000, 10'b1111111111, 10'b1111101100, 10'b1111110000, 10'b0000011110, 10'b0000000000, 10'b1111110111, 10'b1111111111, 10'b0000001101, 10'b1111111111, 10'b1111111111, 10'b1111110010, 10'b0000010100, 10'b0000000000, 10'b0000001001, 10'b1111111110, 10'b0000001010, 10'b0000000000, 10'b0000000000, 10'b0000001111, 10'b1111110011, 10'b1111111101, 10'b0000001010, 10'b1111111001}, 
{10'b1111111110, 10'b1111101100, 10'b0000100110, 10'b1111111011, 10'b0000001100, 10'b1111101101, 10'b0000000000, 10'b0000000010, 10'b1111100001, 10'b1111111111, 10'b1111111000, 10'b0000000011, 10'b1111101011, 10'b0000001000, 10'b0000001100, 10'b0000000111, 10'b0000000101, 10'b1111111101, 10'b1111010010, 10'b1111111111, 10'b1111111100, 10'b0000001000, 10'b1111111000, 10'b1111111111, 10'b0000001100, 10'b1111111101, 10'b1111111111, 10'b0000011000, 10'b1111100110, 10'b1111101101, 10'b0000010110, 10'b0000000010}, 
{10'b0000011011, 10'b0000001100, 10'b0000000000, 10'b1111110101, 10'b1111111010, 10'b1111111111, 10'b0000000000, 10'b1111111011, 10'b1111111000, 10'b1111111000, 10'b0000000000, 10'b0000001010, 10'b0000000000, 10'b0000000011, 10'b1111111101, 10'b0000000000, 10'b1111110110, 10'b0000000000, 10'b1111111110, 10'b1111111111, 10'b0000000000, 10'b0000000011, 10'b0000000110, 10'b0000000000, 10'b0000000000, 10'b1111011000, 10'b1111110011, 10'b0000000000, 10'b0000000001, 10'b0000000000, 10'b1111110100, 10'b0000000001}, 
{10'b0000001100, 10'b1110111101, 10'b1111111111, 10'b1111111011, 10'b1111110001, 10'b1111111111, 10'b0000000000, 10'b0000100011, 10'b1111111101, 10'b1111111110, 10'b0000000101, 10'b1111010101, 10'b0000000001, 10'b1111100011, 10'b0000101110, 10'b1111111100, 10'b1111110001, 10'b1111011100, 10'b1111111111, 10'b1111010010, 10'b1111001100, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b0000001111, 10'b1111111111, 10'b1111101100, 10'b1111111011, 10'b1111111110, 10'b0000000000, 10'b1111111101, 10'b1111010011}
};

localparam logic signed [9:0] bias [32] = '{
10'b0000010000,  // 0.5280959606170654
10'b0000011010,  // 0.8414360880851746
10'b0000001100,  // 0.397830605506897
10'b0000001101,  // 0.4105983078479767
10'b1110001010,  // -3.657735586166382
10'b1111100011,  // -0.8977976441383362
10'b0000110110,  // 1.7051936388015747
10'b1111010111,  // -1.2765135765075684
10'b1111101101,  // -0.5837795734405518
10'b0001010110,  // 2.699671983718872
10'b0000000110,  // 0.2170683741569519
10'b0000011100,  // 0.8814588785171509
10'b1110101011,  // -2.634300947189331
10'b1111000011,  // -1.877297282218933
10'b0000110101,  // 1.6625694036483765
10'b0001010111,  // 2.7459704875946045
10'b1111110000,  // -0.47838035225868225
10'b0000110110,  // 1.6984987258911133
10'b0000011011,  // 0.8548859357833862
10'b0000100000,  // 1.0045719146728516
10'b0000101101,  // 1.4197649955749512
10'b0000011010,  // 0.832463800907135
10'b0000010001,  // 0.5434179306030273
10'b0000011101,  // 0.9277304410934448
10'b1111110101,  // -0.3426123857498169
10'b1111101110,  // -0.5587119460105896
10'b1111101100,  // -0.6208624839782715
10'b1111010111,  // -1.2802538871765137
10'b0000000001,  // 0.05940237268805504
10'b1111100101,  // -0.8213341236114502
10'b0000011100,  // 0.8783953189849854
10'b1111100001   // -0.949700653553009
};
endpackage