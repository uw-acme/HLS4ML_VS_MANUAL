// Width: 16
// NFRAC: 10
package dense_2_16_10;

localparam logic signed [15:0] weights [64][32] = '{ 
{16'b0000000100010011, 16'b0000000000001000, 16'b1111111100111101, 16'b1111111111101010, 16'b0000000100001011, 16'b0000000000000000, 16'b1111111101101100, 16'b1111111111111111, 16'b1111111011100111, 16'b0000000001010001, 16'b0000000000000000, 16'b1111111111111010, 16'b1111111111111111, 16'b1111111100110011, 16'b1111111111001100, 16'b1111111011110011, 16'b0000000000000000, 16'b1111111111110010, 16'b1111111100111100, 16'b1111111101011101, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111110111, 16'b1111111111111101, 16'b0000000000000000, 16'b0000000001100110, 16'b0000000110001011, 16'b0000000010110011, 16'b1111111111111111, 16'b0000000000110011, 16'b1111111001011100, 16'b0000000000000000}, 
{16'b1111111110011001, 16'b1111111101100001, 16'b1111111101110010, 16'b1111111111000111, 16'b1111111111111010, 16'b0000000000101100, 16'b1111111100011011, 16'b0000000000000101, 16'b0000000000000100, 16'b1111111110111111, 16'b0000000010011111, 16'b1111111111010011, 16'b1111111111000011, 16'b1111111100100001, 16'b0000000000000111, 16'b1111111111001110, 16'b0000000000001100, 16'b1111111100111000, 16'b0000000010101111, 16'b0000000011101011, 16'b1111111111011111, 16'b1111111111111010, 16'b1111111111111111, 16'b0000000000011000, 16'b1111111110110111, 16'b0000000100011001, 16'b0000000011111101, 16'b0000000000001000, 16'b0000000000011101, 16'b1111111000001101, 16'b0000000000000111, 16'b0000000000000000}, 
{16'b0000000001001010, 16'b1111111110001010, 16'b1111111101111011, 16'b1111111111010101, 16'b1111111110110000, 16'b1111111110101000, 16'b1111111101000010, 16'b0000000000000100, 16'b1111111101110101, 16'b0000000000001001, 16'b0000000000000010, 16'b1111111110101101, 16'b0000000001011100, 16'b1111111110111101, 16'b1111111111111110, 16'b1111111111011010, 16'b0000000000000101, 16'b0000000001100001, 16'b0000000000111100, 16'b0000000011101011, 16'b0000000000101010, 16'b1111111110101001, 16'b0000000000000000, 16'b0000000000100011, 16'b1111111111101101, 16'b0000000011010110, 16'b0000000010011000, 16'b0000000001100011, 16'b1111111111111111, 16'b1111111101100100, 16'b1111111111110010, 16'b0000000001100101}, 
{16'b0000000010001101, 16'b0000000000010011, 16'b0000000000110110, 16'b1111111111110110, 16'b1111110111110110, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000011100111, 16'b0000000011111000, 16'b1111111111110010, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000101, 16'b1111111111101101, 16'b0000000011011011, 16'b0000000000000000, 16'b1111111111100110, 16'b1111111111111111, 16'b1111111101001011, 16'b1111111111000001, 16'b0000000000110010, 16'b1111111110111111, 16'b1111111111111111, 16'b0000000000000011, 16'b1111111111001100, 16'b0000000001001010, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111100100011, 16'b0000000100111101}, 
{16'b1111110101000101, 16'b1111111111100110, 16'b1111111111111011, 16'b0000000000000101, 16'b1111111111100101, 16'b0000000000000110, 16'b1111111111001101, 16'b1111111101100110, 16'b0000000000110111, 16'b1111111111101011, 16'b1111111111110010, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000011010111, 16'b0000000000000000, 16'b0000000101010000, 16'b1111111111111111, 16'b0000000011011111, 16'b1111111001100110, 16'b0000000000000000, 16'b1111111110001101, 16'b0000000010101100, 16'b0000000100001000, 16'b0000000000000000, 16'b0000000000101110, 16'b0000000010100110, 16'b0000000011110100, 16'b0000000000010001, 16'b1111111111111011, 16'b1111111111111111, 16'b1111111111110001, 16'b0000000011100111}, 
{16'b0000000000111011, 16'b1111111111111111, 16'b0000000010011000, 16'b1111110101100111, 16'b1111101001111101, 16'b1111111010011001, 16'b0000000101101010, 16'b1111110110000010, 16'b1111111111111111, 16'b1111110101001010, 16'b1111110111111110, 16'b1111111010100010, 16'b0000000101101001, 16'b1111111111111111, 16'b1111111111110000, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111101111000, 16'b1111111111111111, 16'b1111111000001011, 16'b0000000000000000, 16'b0000000010111110, 16'b1111111111111111, 16'b0000000000010110, 16'b0000000100010010, 16'b0000000000110100, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000011010010, 16'b1111111111011101, 16'b0000000011001101}, 
{16'b1111111111011011, 16'b1111111101011110, 16'b1111111100001000, 16'b1111111111001111, 16'b1111111011011000, 16'b0000000001000011, 16'b1111111101000111, 16'b1111111101101110, 16'b1111111001010111, 16'b0000000000110001, 16'b1111111111111010, 16'b1111111101011101, 16'b0000000001111001, 16'b1111111111110101, 16'b1111111111010101, 16'b1111110111001001, 16'b1111111111111111, 16'b0000000001010110, 16'b0000000011000100, 16'b1111111101011001, 16'b1111111101100110, 16'b1111111110111111, 16'b1111111111111110, 16'b0000000000011100, 16'b1111111111010001, 16'b1111110101101000, 16'b1111111011110000, 16'b1111111111010001, 16'b0000000000000101, 16'b1111111111101010, 16'b0000000000011111, 16'b1111111111111111}, 
{16'b1111111101100010, 16'b1111111110100011, 16'b1111111110101110, 16'b1111111100001101, 16'b1111111110001001, 16'b1111111111111111, 16'b0000000001101010, 16'b1111111110101111, 16'b0000000011001101, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000011100000, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111110110111, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000101101, 16'b1111111101000111, 16'b0000000000001110, 16'b1111111111111111, 16'b1111111110110110, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111}, 
{16'b1111111000010111, 16'b1111111111000101, 16'b1111111001111010, 16'b0000000001111101, 16'b0000000111110010, 16'b1111111111111111, 16'b1111111111100010, 16'b0000000011110100, 16'b1111111000111110, 16'b1111111111010000, 16'b0000000000000000, 16'b1111111100110001, 16'b1111111111111111, 16'b0000000001001101, 16'b1111111100111100, 16'b0000001100000100, 16'b1111111111110111, 16'b0000000000101111, 16'b0000000011010100, 16'b0000000011111010, 16'b0000000000000000, 16'b1111111010101000, 16'b0000000000000000, 16'b0000000110100101, 16'b1111111101000110, 16'b0000001011001010, 16'b1111111101100111, 16'b1111111100101111, 16'b1111111000011100, 16'b1111111000100100, 16'b0000000000000000, 16'b0000000000110110}, 
{16'b0000000000000000, 16'b1111111111110000, 16'b1111111110110100, 16'b0000000000000000, 16'b0000000100111011, 16'b1111111111101011, 16'b1111111110111110, 16'b0000000001011110, 16'b0000000001100111, 16'b0000000000000011, 16'b1111111111110111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111110001011, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111010, 16'b0000000000000010, 16'b0000000001010110, 16'b0000000000010011, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000111, 16'b0000000000100111, 16'b1111111101111000, 16'b0000000001000101, 16'b0000000011111110, 16'b1111111111111111, 16'b0000000000000110, 16'b0000000000110010, 16'b0000000001000111}, 
{16'b0000000001100010, 16'b0000000000000000, 16'b1111111110010110, 16'b1111111011111111, 16'b1111110011010010, 16'b0000000010001000, 16'b0000000000000000, 16'b1111110010110000, 16'b0000000000100101, 16'b1111111111111111, 16'b0000000000000011, 16'b1111111111111110, 16'b0000000000001010, 16'b0000000000000000, 16'b1111111111101100, 16'b1111111001111001, 16'b1111111111111111, 16'b0000000011100001, 16'b0000000010000001, 16'b0000000011000011, 16'b1111111000111101, 16'b1111111010010011, 16'b0000000001111010, 16'b1111111111011100, 16'b1111111111010000, 16'b0000000101101111, 16'b1111111110011101, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000011011000, 16'b1111111111111111, 16'b0000000000000110}, 
{16'b1111111100110101, 16'b1111111000000111, 16'b0000000000000000, 16'b1111111111111101, 16'b0000000101010100, 16'b1111111011101100, 16'b1111111100011101, 16'b0000000001110110, 16'b1111111111111111, 16'b0000000010011000, 16'b0000000001001011, 16'b1111111110110010, 16'b0000000000000000, 16'b0000000000001110, 16'b1111111111101010, 16'b1111111011111100, 16'b0000000010110011, 16'b0000000000011101, 16'b0000000100110000, 16'b0000000001011000, 16'b0000000000000000, 16'b1111111111011001, 16'b0000000010000001, 16'b1111111110100111, 16'b1111111011000100, 16'b1111111111111001, 16'b0000000010111101, 16'b1111111111111111, 16'b0000000000001000, 16'b1111111110011111, 16'b0000000010001100, 16'b0000000100011010}, 
{16'b0000000000001111, 16'b0000000000000000, 16'b0000000011100000, 16'b0000000000001000, 16'b1111111111010110, 16'b0000000010111000, 16'b0000000001011110, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111101110000, 16'b1111111111001000, 16'b1111111101010100, 16'b1111111111111111, 16'b0000000000110011, 16'b1111111110111001, 16'b0000001101011111, 16'b0000000000000000, 16'b1111111110011111, 16'b1111111100111110, 16'b1111111111110010, 16'b0000000011001011, 16'b0000000010000011, 16'b0000000000000000, 16'b1111111111111101, 16'b0000000011100000, 16'b0000000100010010, 16'b0000000111111011, 16'b0000000000001010, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111110011, 16'b1111111110110110}, 
{16'b1111111101100000, 16'b0000000000110001, 16'b0000000000101000, 16'b1111111100000010, 16'b1111111011101100, 16'b0000000111100000, 16'b0000000000110010, 16'b0000000000000000, 16'b1111111101011011, 16'b1111111110100101, 16'b0000000010000100, 16'b0000000001001000, 16'b0000000000000000, 16'b1111111110101111, 16'b0000000100100100, 16'b1111111111111111, 16'b1111111111110010, 16'b0000000000000000, 16'b0000000000001101, 16'b1111111111010000, 16'b0000000001010000, 16'b0000000000010000, 16'b0000000001110100, 16'b1111111111111111, 16'b0000000000000011, 16'b0000001010100001, 16'b1111111111000110, 16'b1111111111101000, 16'b1111111111111111, 16'b1111111110010000, 16'b1111111111010110, 16'b0000000010110100}, 
{16'b0000000000111100, 16'b0000000001001011, 16'b0000000101001110, 16'b1111111111010111, 16'b0000000001100111, 16'b0000000101100111, 16'b0000000000000000, 16'b1111111111100001, 16'b0000000001111000, 16'b1111111110001011, 16'b1111111111111111, 16'b1111111110000101, 16'b0000000000000000, 16'b0000000110010010, 16'b1111111111101101, 16'b0000000000000001, 16'b0000000011110001, 16'b0000000000000000, 16'b0000000000000011, 16'b1111111010111111, 16'b1111111100000100, 16'b1111111111011011, 16'b1111111111111111, 16'b1111111101101010, 16'b1111111111011011, 16'b1111111110101011, 16'b1111111100110110, 16'b1111111100100110, 16'b0000000000011110, 16'b0000000001110010, 16'b1111111001101001, 16'b0000000000000011}, 
{16'b1111111011001110, 16'b0000000000000000, 16'b1111111111110000, 16'b1111111111001101, 16'b1111111111111111, 16'b0000000010001000, 16'b1111111110110000, 16'b0000000100010101, 16'b1111111010001100, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111100, 16'b1111111110100011, 16'b0000000001010001, 16'b0000000010111011, 16'b1111111111110110, 16'b1111111011111110, 16'b1111111111000011, 16'b0000000001110010, 16'b0000000001000000, 16'b0000000000000000, 16'b0000000000000011, 16'b0000000001010011, 16'b1111111100001010, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000011, 16'b0000000000000000, 16'b1111111101111111}, 
{16'b1111111010100111, 16'b1111111111111010, 16'b1111111111111100, 16'b1111111111101110, 16'b1111111111111011, 16'b0000000001101100, 16'b0000000000000110, 16'b0000000000100011, 16'b0000000000100111, 16'b0000000001000000, 16'b0000000001010000, 16'b0000000010100101, 16'b0000000000011011, 16'b1111111110011100, 16'b0000000000000000, 16'b0000000110000110, 16'b0000000000000000, 16'b0000000000000001, 16'b1111111111111101, 16'b0000000001110000, 16'b0000000010010001, 16'b0000000000011111, 16'b0000000000101010, 16'b1111111111100001, 16'b1111111111011111, 16'b0000000000011011, 16'b1111111110111011, 16'b1111111101111110, 16'b0000000011010110, 16'b1111111111100000, 16'b0000000000100000, 16'b1111111100111111}, 
{16'b0000000000000000, 16'b1111111111111111, 16'b0000000000100110, 16'b0000000000000000, 16'b0000001110100000, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000001110000, 16'b1111111110110011, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000001, 16'b0000000010000100, 16'b0000000000000000, 16'b1111111101101011, 16'b1111111111111111, 16'b1111111110111011, 16'b0000000101001111, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000001000101, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000101010}, 
{16'b1111111111111100, 16'b0000000000011101, 16'b1111111111111111, 16'b0000000000110001, 16'b1111111111010010, 16'b1111111110000101, 16'b1111111111000000, 16'b0000000100011100, 16'b0000000000000000, 16'b0000000001100011, 16'b1111111111110100, 16'b0000000001000010, 16'b1111111111011110, 16'b1111111101011110, 16'b1111111100111100, 16'b0000000000001101, 16'b1111111111111111, 16'b1111111111011100, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000001001101, 16'b0000000000100100, 16'b1111111101111111, 16'b0000000001110010, 16'b1111111101010111, 16'b0000000000000010, 16'b0000000000000000, 16'b1111111101010100, 16'b0000000000000000, 16'b0000000000101110, 16'b1111111111100000}, 
{16'b1111111111110100, 16'b1111111110011010, 16'b0000000000000000, 16'b1111111111000010, 16'b0000000011011101, 16'b1111111111111111, 16'b1111111111101010, 16'b0000000001101101, 16'b1111111001101111, 16'b0000000000000000, 16'b1111111111011000, 16'b1111111111111101, 16'b0000000101100111, 16'b0000000011101010, 16'b1111111110011010, 16'b1111111111101010, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111101110100, 16'b1111111110000110, 16'b0000000010000110, 16'b0000000000000000, 16'b1111111101110011, 16'b0000000000011001, 16'b1111111110101101, 16'b1111111111011101, 16'b0000000010001011, 16'b0000000000000000, 16'b1111111100000010}, 
{16'b0000001010001001, 16'b0000000101011110, 16'b1111111100000000, 16'b0000000000000011, 16'b1111111010011101, 16'b0000000000000000, 16'b0000000011100100, 16'b0000000000011111, 16'b0000000011100101, 16'b1111111111111111, 16'b1111111101100001, 16'b1111111110101111, 16'b0000000010010001, 16'b0000000000011100, 16'b1111111110011011, 16'b0000000010000110, 16'b0000001000100100, 16'b1111111101111010, 16'b1111111011010000, 16'b0000000000000000, 16'b1111111111100010, 16'b1111111101001011, 16'b1111111111110011, 16'b1111111111111110, 16'b0000000001011000, 16'b1111111010001110, 16'b0000000001011011, 16'b1111111111111110, 16'b0000000000000000, 16'b0000000001101111, 16'b1111111111100010, 16'b0000000000111101}, 
{16'b1111111110100001, 16'b1111111100111011, 16'b1111111111011010, 16'b1111111101010100, 16'b1111111111101110, 16'b0000000000110010, 16'b0000000000000000, 16'b1111111111110100, 16'b0000000000100110, 16'b1111111111111100, 16'b0000000000000000, 16'b1111111100100001, 16'b0000000001101000, 16'b0000000001010010, 16'b1111111110010111, 16'b0000000111000110, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111011, 16'b0000000000000000, 16'b0000000101000011, 16'b1111111000011110, 16'b1111111110010001, 16'b1111111111000110, 16'b1111111111101100, 16'b0000000011001001, 16'b1111111111001010, 16'b0000000000010010, 16'b0000000111101111, 16'b1111110111110011, 16'b1111111010001000, 16'b0000000000010110}, 
{16'b0000000000010001, 16'b1111111111000011, 16'b1111111111111111, 16'b0000000000000000, 16'b1111110100011111, 16'b1111110110010011, 16'b0000000000000001, 16'b1111111111111111, 16'b1111111011110000, 16'b0000000000011001, 16'b0000000000000000, 16'b1111111111100011, 16'b0000000000000000, 16'b1111111111000100, 16'b1111111111001010, 16'b1111111110111001, 16'b1111111101101001, 16'b0000000100100001, 16'b0000000000000000, 16'b0000000000101111, 16'b1111111111111111, 16'b1111111110110111, 16'b0000000000000000, 16'b1111111110100111, 16'b0000000011100000, 16'b1111110110000010, 16'b0000000011100001, 16'b1111111111111111, 16'b1111111111111011, 16'b0000000011001100, 16'b1111111111111111, 16'b0000000011110001}, 
{16'b1111111111111111, 16'b0000000000000101, 16'b1111111111010011, 16'b0000000001001100, 16'b0000000000111000, 16'b1111111010100001, 16'b0000000000000000, 16'b0000000001000001, 16'b0000001001010001, 16'b1111111111110110, 16'b0000000000000000, 16'b0000000000111001, 16'b0000000101101111, 16'b1111111111011111, 16'b0000000000001110, 16'b0000000001100111, 16'b1111111111111111, 16'b0000000000011100, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111011100111, 16'b0000000000100111, 16'b0000000001000111, 16'b0000000000010111, 16'b1111111111111111, 16'b0000000011011111, 16'b0000000000000100, 16'b0000000010000001, 16'b1111111001010100, 16'b0000000001101001, 16'b0000000110010101, 16'b0000000000000101}, 
{16'b1111111010011000, 16'b0000000011011000, 16'b1111111011110101, 16'b0000000001111101, 16'b1111111110010100, 16'b0000000000000000, 16'b0000000111111101, 16'b1111111100010001, 16'b1111111011010101, 16'b0000000010101111, 16'b1111111100011011, 16'b1111111111100111, 16'b1111111111111111, 16'b0000000101100000, 16'b1111111111111110, 16'b1111111011001011, 16'b1111111111111111, 16'b0000000111000011, 16'b1111111000011101, 16'b1111111111100111, 16'b0000000101000100, 16'b1111111010001100, 16'b0000000000110110, 16'b1111111111110000, 16'b0000000100010101, 16'b1111110111110111, 16'b1111111010001100, 16'b1111111100110111, 16'b1111111111111111, 16'b0000000001101010, 16'b0000000000011001, 16'b0000000010110110}, 
{16'b1111111110100011, 16'b0000000000110101, 16'b1111111111111111, 16'b0000000010011001, 16'b1111111111011001, 16'b0000000011101000, 16'b0000000000000010, 16'b1111111111110100, 16'b1111111111111101, 16'b0000000000000001, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111110, 16'b0000001000010100, 16'b0000000000001100, 16'b0000000011000001, 16'b0000000000000000, 16'b1111111100100111, 16'b1111111110110001, 16'b1111111111111111, 16'b1111111111101111, 16'b0000000000101011, 16'b1111111111111111, 16'b1111111101000010, 16'b1111111111111111, 16'b0000000100101110, 16'b0000000100111101, 16'b1111111111111111, 16'b1111111111101111, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111110011101}, 
{16'b1111111110101101, 16'b0000000000000000, 16'b0000000100010111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111110001011, 16'b0000000000000000, 16'b1111110010001011, 16'b0000000011011100, 16'b0000000000001110, 16'b0000000000011011, 16'b1111111010001111, 16'b0000000000000011, 16'b1111111101110011, 16'b1111111111011110, 16'b0000000000000000, 16'b0000000000010100, 16'b0000000000000000, 16'b0000000001110011, 16'b0000000000000000, 16'b1111111111110110, 16'b0000000101010001, 16'b0000000110000001, 16'b1111111100011101, 16'b1111111101101110, 16'b0000000011111111, 16'b1111111011000111, 16'b0000000000011110, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000010111100}, 
{16'b1111111110001011, 16'b1111111111111111, 16'b1111111100001011, 16'b1111111100110001, 16'b1111111111110001, 16'b1111111101110101, 16'b0000000000000000, 16'b0000000001011101, 16'b1111111100001010, 16'b1111111110101010, 16'b1111111111001101, 16'b0000000000000000, 16'b0000000000011100, 16'b1111111111110101, 16'b1111111111000001, 16'b0000000001100001, 16'b0000000011100100, 16'b0000000010000110, 16'b1111111101111010, 16'b0000000000110001, 16'b1111111111110011, 16'b1111111111100010, 16'b0000000000010111, 16'b0000000000010000, 16'b1111111110111000, 16'b0000000001011011, 16'b1111111110100011, 16'b0000000000111101, 16'b1111111111111111, 16'b1111111011010001, 16'b1111111111100101, 16'b0000000011100110}, 
{16'b1111111111100100, 16'b1111111110101011, 16'b0000000001001110, 16'b0000000100000011, 16'b0000000001010110, 16'b0000000001010100, 16'b0000000000101111, 16'b1111111100110001, 16'b1111111100101101, 16'b0000000001000110, 16'b0000000000001100, 16'b0000000000101100, 16'b0000000000010110, 16'b0000000000000101, 16'b0000000011010010, 16'b0000000000000111, 16'b1111111111001000, 16'b0000000001101001, 16'b1111111111100001, 16'b1111111111011011, 16'b0000000001110000, 16'b1111111110000001, 16'b1111111111100100, 16'b0000000010000010, 16'b0000000000010110, 16'b1111111110010010, 16'b1111111100110101, 16'b1111111111110011, 16'b1111111011100010, 16'b0000000000111101, 16'b0000000001101000, 16'b0000000000000001}, 
{16'b1111111111110010, 16'b1111111111101011, 16'b1111111111110011, 16'b1111111111011100, 16'b1111111101111001, 16'b1111111101110000, 16'b0000000001000000, 16'b0000000000001000, 16'b1111111101000101, 16'b0000000010101011, 16'b1111111111101010, 16'b1111111111111111, 16'b1111111110001111, 16'b0000000000000101, 16'b0000000000011110, 16'b1111111111001010, 16'b1111111111101111, 16'b1111111111010101, 16'b1111111110101101, 16'b0000000000000000, 16'b1111111101110000, 16'b0000000001101000, 16'b1111111100100111, 16'b0000000000000101, 16'b0000000000101010, 16'b0000000001111110, 16'b0000000000011011, 16'b0000000000000110, 16'b0000000100101011, 16'b0000000000110100, 16'b0000000000000000, 16'b0000000001010101}, 
{16'b1111111111101100, 16'b0000000100000010, 16'b1111111111111111, 16'b1111111111011110, 16'b1111111100100101, 16'b1111111110110011, 16'b0000000110100101, 16'b1111110100111110, 16'b1111111010011010, 16'b1111111100110011, 16'b1111111100011111, 16'b1111111011111100, 16'b1111111111111111, 16'b0000000111101111, 16'b1111111111100101, 16'b0000000000000000, 16'b1111111100100111, 16'b0000000111001000, 16'b1111111001011001, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111010100111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000111001, 16'b1111111111000101, 16'b1111111101101000, 16'b1111111111111111, 16'b0000000010110010, 16'b0000000000000011, 16'b1111111110101101, 16'b0000000000000000}, 
{16'b0000000101111000, 16'b1111111110001101, 16'b0000000010000111, 16'b1111111111011110, 16'b0000000001001110, 16'b1111111111111100, 16'b1111111111111101, 16'b1111111110100000, 16'b0000000000000000, 16'b0000000001011110, 16'b1111111111111111, 16'b1111111111000011, 16'b1111111111111111, 16'b0000000011101010, 16'b0000000000010011, 16'b0000000000101001, 16'b0000000000011000, 16'b1111111111100111, 16'b0000000000010100, 16'b0000000000000000, 16'b1111111111110110, 16'b1111111111111111, 16'b1111111011000111, 16'b1111111111111111, 16'b0000000000111011, 16'b1111111110001000, 16'b1111111101110101, 16'b1111111111111111, 16'b1111111111111111, 16'b0000001000111011, 16'b1111111011011011, 16'b1111111110001001}, 
{16'b1111111111010010, 16'b1111111110010110, 16'b1111111110111101, 16'b0000000000100101, 16'b0000000010001110, 16'b1111111101111011, 16'b1111111111111110, 16'b1111111100011110, 16'b0000000000111110, 16'b0000000010001011, 16'b1111111100100101, 16'b1111111011111101, 16'b0000000000011000, 16'b1111110101000100, 16'b1111111110110010, 16'b1111111110000001, 16'b1111111100110101, 16'b1111111111111111, 16'b0000000010001001, 16'b0000000000000000, 16'b1111111111010001, 16'b1111111111010010, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111000011, 16'b1111110011111011, 16'b1111110111000111, 16'b1111111011101000, 16'b0000000000111001, 16'b0000000011010011, 16'b1111111111111111, 16'b0000000011110110}, 
{16'b1111111110100001, 16'b1111111100100100, 16'b0000000010100111, 16'b0000000001001100, 16'b0000000000101100, 16'b1111111110100001, 16'b1111111111011110, 16'b0000000001100100, 16'b0000001000100111, 16'b1111111101010000, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000001111000, 16'b1111111111000111, 16'b1111111111101101, 16'b1111111111101110, 16'b1111111110011001, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000011101000, 16'b1111111101110111, 16'b1111111111111100, 16'b0000000010000011, 16'b1111111111110101, 16'b0000000000000000, 16'b0000001000011010, 16'b0000000101001100, 16'b0000000000000011, 16'b0000000000000000, 16'b1111111001010001, 16'b1111111110111010, 16'b1111111111111111}, 
{16'b0000000000001111, 16'b0000000000110001, 16'b1111111111110001, 16'b0000000000000000, 16'b0000000011101100, 16'b1111111000010001, 16'b0000000000000000, 16'b1111111110011110, 16'b0000000010111110, 16'b0000000000000000, 16'b1111111111101101, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000101, 16'b1111111110010001, 16'b0000000100001001, 16'b1111111111111010, 16'b1111111111110000, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000001101, 16'b1111111010111011, 16'b0000000000110100, 16'b0000000010111011, 16'b1111111111111100, 16'b0000000001100000, 16'b1111111111111111, 16'b0000000001001100}, 
{16'b1111111100110001, 16'b0000000000001001, 16'b1111111000010010, 16'b0000000000000111, 16'b1111111111001100, 16'b1111111111010111, 16'b1111111111111110, 16'b1111111110100010, 16'b1111111111011011, 16'b1111111110111101, 16'b0000000000110000, 16'b0000000000011011, 16'b1111111101001010, 16'b0000000000000000, 16'b1111111111111110, 16'b1111111111110111, 16'b0000000001001000, 16'b1111111111101011, 16'b1111111111100011, 16'b1111111111100010, 16'b1111111111111111, 16'b0000000100010101, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111110110, 16'b0000000101000100, 16'b0000000011000001, 16'b0000000000100010, 16'b1111111110011101, 16'b1111111111110101, 16'b0000000001000010, 16'b0000000000111010}, 
{16'b0000000000100010, 16'b0000000000101000, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111000100000, 16'b0000000000101100, 16'b0000000000011001, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111101010010, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111101011011, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111010010011, 16'b0000000000001001, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000010000100, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000111010010, 16'b0000000101011100, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111100010000, 16'b0000000000000000, 16'b1111111111111111}, 
{16'b0000000001001101, 16'b0000000000110110, 16'b0000000100000011, 16'b1111111100000001, 16'b0000000010000111, 16'b0000000001111001, 16'b0000000000000110, 16'b0000000011000100, 16'b0000000000001100, 16'b1111111111110011, 16'b0000000000100110, 16'b0000000000000101, 16'b1111111111111111, 16'b0000000001111011, 16'b1111111111111010, 16'b1111111111010111, 16'b0000000000000000, 16'b0000000000100000, 16'b1111111111001110, 16'b0000000001100101, 16'b0000000000100001, 16'b1111110110101101, 16'b1111111110001010, 16'b0000000001011101, 16'b1111111111111111, 16'b1111110111111010, 16'b1111111101111110, 16'b1111111111101000, 16'b1111111111111111, 16'b1111111111000101, 16'b0000000000000000, 16'b1111111111010111}, 
{16'b0000000000000001, 16'b1111111111111111, 16'b1111111110100010, 16'b1111111101010011, 16'b0000000000101010, 16'b0000000000000000, 16'b0000000001100001, 16'b1111111111111010, 16'b0000000011111111, 16'b1111111111111011, 16'b0000000000000000, 16'b1111111010100000, 16'b1111111111111111, 16'b0000000010000000, 16'b1111111111111111, 16'b1111111011110101, 16'b0000000000000000, 16'b1111111111110100, 16'b0000000100001101, 16'b1111111111111111, 16'b1111111001000000, 16'b1111111111111111, 16'b0000000100001000, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000010001110, 16'b1111111110011111, 16'b0000000001000110, 16'b0000000000000000, 16'b1111111100110001, 16'b0000000000000000, 16'b0000000000000010}, 
{16'b1111111100100010, 16'b0000000000000001, 16'b0000000000000000, 16'b1111111111111001, 16'b0000000111111011, 16'b1111111110000000, 16'b1111111111111010, 16'b1111111111111000, 16'b1111111111010010, 16'b1111111111001100, 16'b0000000001000010, 16'b0000000010001000, 16'b1111111111011010, 16'b0000000011111111, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111011011101, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111110101110, 16'b0000000000000010, 16'b0000000000100110, 16'b0000000000001101, 16'b1111111111110110, 16'b1111111111001011, 16'b1111111100110000, 16'b1111111011010001, 16'b0000000000000000, 16'b1111111110001100, 16'b0000000000101000, 16'b1111111111111111, 16'b0000000001001101}, 
{16'b1111111001011000, 16'b1111111101011111, 16'b1111111101100000, 16'b0000000000000000, 16'b0000001001001000, 16'b1111111100011100, 16'b0000000000000000, 16'b1111111111001000, 16'b1111111001011100, 16'b0000000010001101, 16'b1111111111111111, 16'b0000001001000100, 16'b0000000000000000, 16'b1111111111001111, 16'b1111111111111111, 16'b0000000000100000, 16'b1111111111101100, 16'b0000000000000000, 16'b1111111111010000, 16'b0000000111111011, 16'b0000000000100111, 16'b1111111111010101, 16'b0000000001110000, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111110011100, 16'b1111111111010000, 16'b1111111000100000, 16'b1111111101101100, 16'b1111111111111111, 16'b1111111111111110, 16'b1111111111000011}, 
{16'b0000000011100111, 16'b1111110011001101, 16'b1111110100011010, 16'b1111111101010001, 16'b0000001010101101, 16'b1111111111111111, 16'b1111111010011101, 16'b0000000100001111, 16'b0000000000111100, 16'b0000000000000000, 16'b0000000011010101, 16'b1111111011101010, 16'b0000000000000000, 16'b0000000000000100, 16'b1111111111011111, 16'b0000000000010010, 16'b1111111110010101, 16'b1111110001010000, 16'b0000000010101011, 16'b0000000101100001, 16'b0000000100001111, 16'b0000000000000010, 16'b0000000000011101, 16'b1111111001100011, 16'b1111110101111000, 16'b1111111111111010, 16'b1111111011001101, 16'b1111111000101011, 16'b1111111100111000, 16'b1111110001111101, 16'b0000000110101101, 16'b0000000110110111}, 
{16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000010, 16'b0000000000000000, 16'b0000000100001001, 16'b1111111101000000, 16'b0000000000010010, 16'b0000000001001010, 16'b1111111010011010, 16'b0000000000100101, 16'b1111111111111011, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000011110101, 16'b0000000000110101, 16'b0000000000010110, 16'b0000000000111111, 16'b0000000101010101, 16'b1111111100100000, 16'b0000000000000000, 16'b1111111101010111, 16'b1111111111111111, 16'b0000000101000010, 16'b0000000000001000, 16'b1111111111111101, 16'b1111110111000001, 16'b1111111111110110, 16'b1111111101100001, 16'b1111111111000001, 16'b0000000000000011, 16'b0000000010001010, 16'b0000000001101010}, 
{16'b1111111111010011, 16'b0000000010001001, 16'b1111111011001000, 16'b0000000000010101, 16'b0000000011000110, 16'b1111111111010111, 16'b1111111111111011, 16'b0000000010100111, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111110111101, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111011100, 16'b1111111110000011, 16'b1111111110111100, 16'b1111111111000110, 16'b1111111110111111, 16'b1111111110001111, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111010010, 16'b1111111110111011, 16'b0000000110010111, 16'b0000000000000000, 16'b1111111010001111, 16'b1111111111110111, 16'b0000000001111110, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000100000000, 16'b1111111111111111}, 
{16'b1111111111111111, 16'b0000000000000100, 16'b1111111111111111, 16'b1111111101100000, 16'b1111110010001111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111001, 16'b1111110110011010, 16'b0000000001010011, 16'b1111111110011011, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111010000101, 16'b1111111111010001, 16'b1111111111111111, 16'b0000000000000001, 16'b0000000000001000, 16'b0000000000100101, 16'b0000000101100001, 16'b1111111110000101, 16'b1111111011001101, 16'b0000000000000000, 16'b1111111011110111, 16'b1111111110011010, 16'b1111111100010011, 16'b1111111111111000, 16'b1111111111110011, 16'b1111111111101101, 16'b1111111000011101, 16'b1111111111011101, 16'b0000000011111000}, 
{16'b0000000001110011, 16'b0000000011100000, 16'b1111111111111101, 16'b0000000010100011, 16'b1111111100101000, 16'b1111111110000000, 16'b0000000001100001, 16'b0000000001000110, 16'b1111111111001111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111010110111, 16'b1111111111111111, 16'b0000000010010011, 16'b1111111110001010, 16'b0000000000100011, 16'b1111111111111110, 16'b1111111111111110, 16'b0000000011010100, 16'b1111111010110001, 16'b0000000100011111, 16'b0000000000110000, 16'b0000000000000000, 16'b0000000011011000, 16'b0000000000000011, 16'b1111111111011011, 16'b1111111001111010, 16'b1111111110001111, 16'b1111111101010001, 16'b0000000010110101}, 
{16'b0000000000000000, 16'b0000000000000111, 16'b1111111010001001, 16'b1111111111111101, 16'b0000000011010011, 16'b1111111101101111, 16'b1111111111110011, 16'b1111111111111111, 16'b0000000000010100, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111100101111, 16'b0000000001100010, 16'b0000000000000110, 16'b0000000000000000, 16'b0000000000100110, 16'b1111111111111111, 16'b1111111101100111, 16'b0000000000010010, 16'b0000000000000000, 16'b1111111111011100, 16'b1111111111101001, 16'b0000000100101111, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111011010100, 16'b1111111010110001, 16'b0000000011110111, 16'b1111111111111110, 16'b1111111111111111, 16'b0000000000011100, 16'b0000000100100001}, 
{16'b1111111010100011, 16'b1111111111111111, 16'b1111111100100110, 16'b0000000000000100, 16'b1111111010010110, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111110111101, 16'b1111110111011110, 16'b1111111111100101, 16'b0000000000000000, 16'b1111111111110111, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111110111, 16'b1111111111001101, 16'b1111111101101000, 16'b1111111110011110, 16'b0000000001000011, 16'b1111111111111101, 16'b1111111111100110, 16'b0000000000000000, 16'b0000000101011000, 16'b1111111111111111, 16'b0000000010011001, 16'b0000000001011101, 16'b1111111101110011, 16'b0000000011011010, 16'b1111111111010001, 16'b0000000000000000, 16'b1111111111111110, 16'b0000001001010100}, 
{16'b1111111010111110, 16'b0000000000011110, 16'b0000000000110011, 16'b1111111111100011, 16'b0000000011111010, 16'b1111111011001010, 16'b1111111111111000, 16'b0000000100001111, 16'b0000000010100011, 16'b0000000000001001, 16'b1111111111111111, 16'b1111111110111001, 16'b1111111110100100, 16'b1111111110111101, 16'b1111111111001101, 16'b0000000001011100, 16'b1111111111111111, 16'b0000000000001000, 16'b0000000010010000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000001111, 16'b0000000100000010, 16'b0000000000101110, 16'b0000000000000110, 16'b1111111110010001, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111110001, 16'b1111111111110011, 16'b1111111111111111, 16'b0000000001000101}, 
{16'b1111111111111111, 16'b0000000000000011, 16'b1111111100100110, 16'b1111111110110011, 16'b0000000100100000, 16'b1111111111111111, 16'b1111111110110000, 16'b0000000011111010, 16'b1111111111001001, 16'b0000000100101010, 16'b0000000001010111, 16'b1111111110000100, 16'b0000000000000000, 16'b0000000000000011, 16'b1111111111110000, 16'b0000000000010101, 16'b1111111110110001, 16'b1111111011110010, 16'b0000000100011100, 16'b0000000010011111, 16'b0000001010001001, 16'b0000000011001101, 16'b0000000011111110, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000111010, 16'b0000000001010001, 16'b1111111001010001, 16'b1111111111111111, 16'b1111111111111010, 16'b1111111111111001}, 
{16'b0000000000000000, 16'b1111111110100110, 16'b1111111110010101, 16'b0000000000000000, 16'b1111111100000110, 16'b0000000000000000, 16'b0000000011000100, 16'b0000000001101111, 16'b0000000000110110, 16'b1111111110011010, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111010100, 16'b0000000011001110, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111011001010, 16'b0000000000000000, 16'b1111111100111010, 16'b1111111111111110, 16'b0000000000000000, 16'b1111111111111011, 16'b0000000000001111, 16'b0000000000010001, 16'b0000000000011100, 16'b0000000010001101, 16'b1111111110111101, 16'b1111111111111000, 16'b1111111000110100, 16'b0000000001010000}, 
{16'b0000000111000100, 16'b1111111111110111, 16'b0000000001000011, 16'b1111111110010100, 16'b1111111110101000, 16'b0000000000100010, 16'b0000000010100100, 16'b0000000000000000, 16'b0000001000011011, 16'b0000000000000000, 16'b1111111111101010, 16'b0000000000010011, 16'b0000000001100000, 16'b1111111111111101, 16'b0000000000110110, 16'b0000000001101001, 16'b1111111111111011, 16'b1111111000111000, 16'b1111111111000110, 16'b1111111111111110, 16'b0000000001110111, 16'b0000000000000001, 16'b1111111111111111, 16'b0000000001110011, 16'b0000000000010010, 16'b1111111011110010, 16'b1111111110010110, 16'b0000000010000111, 16'b1111111111100011, 16'b0000000100001000, 16'b1111111111111110, 16'b1111111101001000}, 
{16'b0000000000001101, 16'b0000000001101000, 16'b1111111111111111, 16'b1111111111011000, 16'b1111111010010110, 16'b1111111111111111, 16'b0000000000101111, 16'b1111111111010000, 16'b0000000010101000, 16'b1111111111011101, 16'b1111111111111111, 16'b1111111111011101, 16'b1111111111111111, 16'b1111111111011010, 16'b0000000000000000, 16'b0000000101000000, 16'b0000000000000000, 16'b1111111111111110, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000100010, 16'b0000000010000000, 16'b0000000000000000, 16'b0000000000000100, 16'b0000000000100001, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000010100, 16'b0000000000000001, 16'b0000000001100011}, 
{16'b1111111011000011, 16'b0000000010000101, 16'b0000000000010010, 16'b1111111110010100, 16'b1111111001100111, 16'b1111111111101101, 16'b0000000001000100, 16'b1111111001101001, 16'b0000001000001011, 16'b0000000001001001, 16'b0000000000010000, 16'b0000000001100000, 16'b0000000000101101, 16'b0000000000000000, 16'b0000000110100001, 16'b1111111110101001, 16'b0000000000000101, 16'b0000000000000000, 16'b1111111111111001, 16'b0000000000000011, 16'b1111111001000101, 16'b0000000000010001, 16'b0000000010011100, 16'b0000000000100110, 16'b0000000000100100, 16'b1111110101011111, 16'b1111111010100010, 16'b1111111100001001, 16'b0000000000000010, 16'b1111111111111110, 16'b0000000101001101, 16'b1111111100101110}, 
{16'b1111111111110010, 16'b1111111100111000, 16'b1111111110010110, 16'b1111111001011101, 16'b1111111011110101, 16'b0000000101011000, 16'b0000000100111101, 16'b1111111101010001, 16'b0000000000101010, 16'b1111111111011000, 16'b1111111110011111, 16'b1111111011111110, 16'b0000000001101001, 16'b1111111011011101, 16'b0000000011000001, 16'b1111111111111111, 16'b0000000101010111, 16'b1111111111111111, 16'b1111111111111000, 16'b1111111101110101, 16'b1111111111010101, 16'b1111111110111101, 16'b1111111011101111, 16'b0000000001010100, 16'b1111111111111111, 16'b1111111111111001, 16'b1111111100010110, 16'b0000000101000010, 16'b0000000100011101, 16'b1111111110100011, 16'b1111110101111010, 16'b0000000010010010}, 
{16'b0000000000000000, 16'b1111111111100101, 16'b1111111111111111, 16'b1111111110011100, 16'b0000000000011101, 16'b0000000000001001, 16'b0000000001000111, 16'b0000000000000101, 16'b0000000001111000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000001100001, 16'b0000000000000001, 16'b0000000000001100, 16'b1111111101111000, 16'b1111111110010001, 16'b0000000000000000, 16'b0000000010111010, 16'b0000000000111010, 16'b0000000010000000, 16'b1111111111101111, 16'b1111111101011100, 16'b1111111111111111, 16'b0000000001001100, 16'b1111111111111111, 16'b0000000000100001, 16'b1111111111111011, 16'b0000000001000101, 16'b0000000000000000, 16'b0000000001010101, 16'b1111111001111011, 16'b1111111111111111}, 
{16'b0000000100111101, 16'b1111111111110110, 16'b0000000010011001, 16'b1111111011000111, 16'b1111111100111010, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000011100, 16'b0000000000000010, 16'b1111111101111111, 16'b0000000000000000, 16'b0000000000000010, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111101111011, 16'b0000000010010010, 16'b1111111111111110, 16'b1111111111100000, 16'b0000000000000000, 16'b0000000001111010, 16'b1111111100110010, 16'b0000000001110110, 16'b0000000010001111, 16'b0000000010000100, 16'b1111111111111111, 16'b0000001000110100, 16'b1111111101100011, 16'b0000000101110100, 16'b1111111111001011, 16'b1111111010001110, 16'b1111111101001110, 16'b0000000010001110}, 
{16'b1111110111010011, 16'b1111111111100100, 16'b1111111101100010, 16'b1111111111111111, 16'b0000000100001011, 16'b1111111101001001, 16'b1111111111000010, 16'b0000000011110011, 16'b0000000001100000, 16'b1111111100001100, 16'b0000000000000000, 16'b1111111111100011, 16'b1111111111110101, 16'b0000000010001100, 16'b1111111100000100, 16'b1111111111110100, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111101111, 16'b0000000000000000, 16'b1111111100111101, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111010101111, 16'b0000000001000111, 16'b0000001001111010, 16'b0000000101100010, 16'b1111111111011011, 16'b1111111101011011, 16'b1111111000110100, 16'b0000000000000000, 16'b1111111111001110}, 
{16'b0000000000010101, 16'b0000000011011010, 16'b0000000000010101, 16'b1111111101100101, 16'b0000000000000100, 16'b1111111111100101, 16'b0000000000000000, 16'b0000000011010101, 16'b0000000011011100, 16'b1111111101110111, 16'b0000000010001111, 16'b0000000000011000, 16'b1111111111111111, 16'b1111111111110001, 16'b1111111101011101, 16'b0000000100000011, 16'b1111111111010100, 16'b1111111010110101, 16'b0000000001110101, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000001110111, 16'b1111111110110011, 16'b1111111111111011, 16'b1111111111001011, 16'b0000000001011010, 16'b1111111101110000, 16'b0000000010001001, 16'b1111111010001011, 16'b0000000001010010, 16'b1111111111111111, 16'b0000000010100000}, 
{16'b1111111111010100, 16'b0000000000000000, 16'b0000000001011011, 16'b0000000000000000, 16'b1111111111000001, 16'b1111111111111101, 16'b0000000001101001, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000101, 16'b0000000000000000, 16'b0000000000010100, 16'b1111111110010011, 16'b0000000000001010, 16'b0000000001110001, 16'b0000000000101111, 16'b0000000001101100, 16'b1111111111111111, 16'b1111111111111110, 16'b0000000010000011, 16'b0000000011111101, 16'b1111111110011011, 16'b0000000000000000, 16'b1111111111111101, 16'b0000000000001011, 16'b1111111000100111, 16'b1111111111111111, 16'b1111111110110111, 16'b1111111111111111, 16'b0000001001000010, 16'b0000000000000000, 16'b1111111100101101}, 
{16'b1111111111100100, 16'b1111111110000101, 16'b1111111111110110, 16'b0000000000000111, 16'b0000000001011100, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111101000, 16'b0000000001001000, 16'b1111111111110111, 16'b0000000000000000, 16'b0000000000100000, 16'b0000000100101110, 16'b1111111110010111, 16'b0000000000001100, 16'b1111110010011011, 16'b1111111111110100, 16'b1111111111000010, 16'b0000000000001000, 16'b1111111111001100, 16'b0000000001011110, 16'b1111111100011010, 16'b0000000001110100, 16'b0000000001101011, 16'b1111111111110010, 16'b1111110100100111, 16'b1111111100010101, 16'b1111111111101001, 16'b1111111111101101, 16'b0000000110001111, 16'b1111111111111010, 16'b0000000010011101}, 
{16'b0000000000110000, 16'b0000000000000000, 16'b0000000010110010, 16'b1111111110001011, 16'b1111111110111001, 16'b0000000011110011, 16'b1111111101011100, 16'b0000000000111010, 16'b1111111011000011, 16'b0000000000001000, 16'b0000000000010001, 16'b1111111110101010, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111100111111, 16'b0000000110111010, 16'b1111111100000011, 16'b1111111111110011, 16'b0000000001111001, 16'b1111111111111111, 16'b0000000001000110, 16'b1111111000010101, 16'b0000000101000000, 16'b1111111111111111, 16'b1111111110000001, 16'b0000000111110000, 16'b0000000010010101, 16'b1111111101011110, 16'b1111111101110110, 16'b1111110111011001, 16'b1111111111110101, 16'b0000000000010000}, 
{16'b1111111111111111, 16'b0000000000000110, 16'b1111111111011100, 16'b1111111011101101, 16'b1111111111111111, 16'b1111111001101110, 16'b0000000000000000, 16'b0000000100110110, 16'b0000000011111010, 16'b0000000000010011, 16'b0000000000000000, 16'b1111111110001111, 16'b0000000101010100, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000110111100, 16'b0000000000000001, 16'b1111111111010111, 16'b1111111111001011, 16'b1111111010110110, 16'b0000000010000110, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000100000, 16'b1111111110110111, 16'b1111111000101000, 16'b0000000100011010, 16'b1111111000111001, 16'b0000000000110100, 16'b1111111110101111, 16'b0000000000000000}, 
{16'b0000000000111110, 16'b0000000010111110, 16'b0000000000001001, 16'b1111111111111100, 16'b1111111000101001, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000011111000, 16'b0000000100011011, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111110, 16'b0000000000000000, 16'b0000000000000010, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000010101110, 16'b1111111110010110, 16'b1111111001000101, 16'b1111111111011110, 16'b1111111110011010, 16'b1111111110011111, 16'b1111111110111001, 16'b1111111111111111, 16'b1111111110111111, 16'b1111111111101001, 16'b1111111111110101, 16'b0000000010010000, 16'b1111111111111111, 16'b0000000111011010}
};

localparam logic signed [15:0] bias [32] = '{
16'b0000010111100101,  // 1.474280834197998
16'b0000001011000100,  // 0.6914801001548767
16'b0000010111000011,  // 1.4406442642211914
16'b0000010110100001,  // 1.408045768737793
16'b0000001111110010,  // 0.9864811301231384
16'b0000001101110100,  // 0.8636202812194824
16'b1111110110001001,  // -0.6153604388237
16'b0000000111101111,  // 0.4839226007461548
16'b0000000111110001,  // 0.4862793982028961
16'b0000000101111100,  // 0.37162142992019653
16'b0000000111010110,  // 0.45989668369293213
16'b0000010100110011,  // 1.2998151779174805
16'b1111101111101111,  // -1.016528844833374
16'b1111111010010111,  // -0.35249894857406616
16'b0000000111001000,  // 0.44582197070121765
16'b1111111110001101,  // -0.1119980737566948
16'b1111111110111011,  // -0.06717441976070404
16'b0000000000000100,  // 0.00487547367811203
16'b0000000011000111,  // 0.1946917623281479
16'b1111110011100001,  // -0.7796769738197327
16'b0000001011101010,  // 0.7287401556968689
16'b0000011011011100,  // 1.714877724647522
16'b1111100110011100,  // -1.5971007347106934
16'b0000000001001011,  // 0.07393483817577362
16'b0000000101001010,  // 0.3225609362125397
16'b0000001101100001,  // 0.8453295230865479
16'b0000001110011000,  // 0.898597240447998
16'b0000000100000100,  // 0.2548799514770508
16'b0000001111100100,  // 0.9735668301582336
16'b0000010010000001,  // 1.1261906623840332
16'b0000000111001010,  // 0.44768181443214417
16'b1111011010000111   // -2.3676068782806396
};
endpackage