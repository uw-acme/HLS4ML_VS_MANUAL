// Width: 16
// NFRAC: 8
package dense_2_16_8;

localparam logic signed [15:0] weights [64][32] = '{ 
{16'b0000000001000100, 16'b0000000000000010, 16'b1111111111001111, 16'b1111111111111010, 16'b0000000001000010, 16'b0000000000000000, 16'b1111111111011011, 16'b1111111111111111, 16'b1111111110111001, 16'b0000000000010100, 16'b0000000000000000, 16'b1111111111111110, 16'b1111111111111111, 16'b1111111111001100, 16'b1111111111110011, 16'b1111111110111100, 16'b0000000000000000, 16'b1111111111111100, 16'b1111111111001111, 16'b1111111111010111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111101, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000011001, 16'b0000000001100010, 16'b0000000000101100, 16'b1111111111111111, 16'b0000000000001100, 16'b1111111110010111, 16'b0000000000000000}, 
{16'b1111111111100110, 16'b1111111111011000, 16'b1111111111011100, 16'b1111111111110001, 16'b1111111111111110, 16'b0000000000001011, 16'b1111111111000110, 16'b0000000000000001, 16'b0000000000000001, 16'b1111111111101111, 16'b0000000000100111, 16'b1111111111110100, 16'b1111111111110000, 16'b1111111111001000, 16'b0000000000000001, 16'b1111111111110011, 16'b0000000000000011, 16'b1111111111001110, 16'b0000000000101011, 16'b0000000000111010, 16'b1111111111110111, 16'b1111111111111110, 16'b1111111111111111, 16'b0000000000000110, 16'b1111111111101101, 16'b0000000001000110, 16'b0000000000111111, 16'b0000000000000010, 16'b0000000000000111, 16'b1111111110000011, 16'b0000000000000001, 16'b0000000000000000}, 
{16'b0000000000010010, 16'b1111111111100010, 16'b1111111111011110, 16'b1111111111110101, 16'b1111111111101100, 16'b1111111111101010, 16'b1111111111010000, 16'b0000000000000001, 16'b1111111111011101, 16'b0000000000000010, 16'b0000000000000000, 16'b1111111111101011, 16'b0000000000010111, 16'b1111111111101111, 16'b1111111111111111, 16'b1111111111110110, 16'b0000000000000001, 16'b0000000000011000, 16'b0000000000001111, 16'b0000000000111010, 16'b0000000000001010, 16'b1111111111101010, 16'b0000000000000000, 16'b0000000000001000, 16'b1111111111111011, 16'b0000000000110101, 16'b0000000000100110, 16'b0000000000011000, 16'b1111111111111111, 16'b1111111111011001, 16'b1111111111111100, 16'b0000000000011001}, 
{16'b0000000000100011, 16'b0000000000000100, 16'b0000000000001101, 16'b1111111111111101, 16'b1111111101111101, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000111001, 16'b0000000000111110, 16'b1111111111111100, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000001, 16'b1111111111111011, 16'b0000000000110110, 16'b0000000000000000, 16'b1111111111111001, 16'b1111111111111111, 16'b1111111111010010, 16'b1111111111110000, 16'b0000000000001100, 16'b1111111111101111, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111110011, 16'b0000000000010010, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111001000, 16'b0000000001001111}, 
{16'b1111111101010001, 16'b1111111111111001, 16'b1111111111111110, 16'b0000000000000001, 16'b1111111111111001, 16'b0000000000000001, 16'b1111111111110011, 16'b1111111111011001, 16'b0000000000001101, 16'b1111111111111010, 16'b1111111111111100, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000110101, 16'b0000000000000000, 16'b0000000001010100, 16'b1111111111111111, 16'b0000000000110111, 16'b1111111110011001, 16'b0000000000000000, 16'b1111111111100011, 16'b0000000000101011, 16'b0000000001000010, 16'b0000000000000000, 16'b0000000000001011, 16'b0000000000101001, 16'b0000000000111101, 16'b0000000000000100, 16'b1111111111111110, 16'b1111111111111111, 16'b1111111111111100, 16'b0000000000111001}, 
{16'b0000000000001110, 16'b1111111111111111, 16'b0000000000100110, 16'b1111111101011001, 16'b1111111010011111, 16'b1111111110100110, 16'b0000000001011010, 16'b1111111101100000, 16'b1111111111111111, 16'b1111111101010010, 16'b1111111101111111, 16'b1111111110101000, 16'b0000000001011010, 16'b1111111111111111, 16'b1111111111111100, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111011110, 16'b1111111111111111, 16'b1111111110000010, 16'b0000000000000000, 16'b0000000000101111, 16'b1111111111111111, 16'b0000000000000101, 16'b0000000001000100, 16'b0000000000001101, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000110100, 16'b1111111111110111, 16'b0000000000110011}, 
{16'b1111111111110110, 16'b1111111111010111, 16'b1111111111000010, 16'b1111111111110011, 16'b1111111110110110, 16'b0000000000010000, 16'b1111111111010001, 16'b1111111111011011, 16'b1111111110010101, 16'b0000000000001100, 16'b1111111111111110, 16'b1111111111010111, 16'b0000000000011110, 16'b1111111111111101, 16'b1111111111110101, 16'b1111111101110010, 16'b1111111111111111, 16'b0000000000010101, 16'b0000000000110001, 16'b1111111111010110, 16'b1111111111011001, 16'b1111111111101111, 16'b1111111111111111, 16'b0000000000000111, 16'b1111111111110100, 16'b1111111101011010, 16'b1111111110111100, 16'b1111111111110100, 16'b0000000000000001, 16'b1111111111111010, 16'b0000000000000111, 16'b1111111111111111}, 
{16'b1111111111011000, 16'b1111111111101000, 16'b1111111111101011, 16'b1111111111000011, 16'b1111111111100010, 16'b1111111111111111, 16'b0000000000011010, 16'b1111111111101011, 16'b0000000000110011, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000111000, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111101101, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000001011, 16'b1111111111010001, 16'b0000000000000011, 16'b1111111111111111, 16'b1111111111101101, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111}, 
{16'b1111111110000101, 16'b1111111111110001, 16'b1111111110011110, 16'b0000000000011111, 16'b0000000001111100, 16'b1111111111111111, 16'b1111111111111000, 16'b0000000000111101, 16'b1111111110001111, 16'b1111111111110100, 16'b0000000000000000, 16'b1111111111001100, 16'b1111111111111111, 16'b0000000000010011, 16'b1111111111001111, 16'b0000000011000001, 16'b1111111111111101, 16'b0000000000001011, 16'b0000000000110101, 16'b0000000000111110, 16'b0000000000000000, 16'b1111111110101010, 16'b0000000000000000, 16'b0000000001101001, 16'b1111111111010001, 16'b0000000010110010, 16'b1111111111011001, 16'b1111111111001011, 16'b1111111110000111, 16'b1111111110001001, 16'b0000000000000000, 16'b0000000000001101}, 
{16'b0000000000000000, 16'b1111111111111100, 16'b1111111111101101, 16'b0000000000000000, 16'b0000000001001110, 16'b1111111111111010, 16'b1111111111101111, 16'b0000000000010111, 16'b0000000000011001, 16'b0000000000000000, 16'b1111111111111101, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111100010, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111110, 16'b0000000000000000, 16'b0000000000010101, 16'b0000000000000100, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000001, 16'b0000000000001001, 16'b1111111111011110, 16'b0000000000010001, 16'b0000000000111111, 16'b1111111111111111, 16'b0000000000000001, 16'b0000000000001100, 16'b0000000000010001}, 
{16'b0000000000011000, 16'b0000000000000000, 16'b1111111111100101, 16'b1111111110111111, 16'b1111111100110100, 16'b0000000000100010, 16'b0000000000000000, 16'b1111111100101100, 16'b0000000000001001, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000010, 16'b0000000000000000, 16'b1111111111111011, 16'b1111111110011110, 16'b1111111111111111, 16'b0000000000111000, 16'b0000000000100000, 16'b0000000000110000, 16'b1111111110001111, 16'b1111111110100100, 16'b0000000000011110, 16'b1111111111110111, 16'b1111111111110100, 16'b0000000001011011, 16'b1111111111100111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000110110, 16'b1111111111111111, 16'b0000000000000001}, 
{16'b1111111111001101, 16'b1111111110000001, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000001010101, 16'b1111111110111011, 16'b1111111111000111, 16'b0000000000011101, 16'b1111111111111111, 16'b0000000000100110, 16'b0000000000010010, 16'b1111111111101100, 16'b0000000000000000, 16'b0000000000000011, 16'b1111111111111010, 16'b1111111110111111, 16'b0000000000101100, 16'b0000000000000111, 16'b0000000001001100, 16'b0000000000010110, 16'b0000000000000000, 16'b1111111111110110, 16'b0000000000100000, 16'b1111111111101001, 16'b1111111110110001, 16'b1111111111111110, 16'b0000000000101111, 16'b1111111111111111, 16'b0000000000000010, 16'b1111111111100111, 16'b0000000000100011, 16'b0000000001000110}, 
{16'b0000000000000011, 16'b0000000000000000, 16'b0000000000111000, 16'b0000000000000010, 16'b1111111111110101, 16'b0000000000101110, 16'b0000000000010111, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111011100, 16'b1111111111110010, 16'b1111111111010101, 16'b1111111111111111, 16'b0000000000001100, 16'b1111111111101110, 16'b0000000011010111, 16'b0000000000000000, 16'b1111111111100111, 16'b1111111111001111, 16'b1111111111111100, 16'b0000000000110010, 16'b0000000000100000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000111000, 16'b0000000001000100, 16'b0000000001111110, 16'b0000000000000010, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111100, 16'b1111111111101101}, 
{16'b1111111111011000, 16'b0000000000001100, 16'b0000000000001010, 16'b1111111111000000, 16'b1111111110111011, 16'b0000000001111000, 16'b0000000000001100, 16'b0000000000000000, 16'b1111111111010110, 16'b1111111111101001, 16'b0000000000100001, 16'b0000000000010010, 16'b0000000000000000, 16'b1111111111101011, 16'b0000000001001001, 16'b1111111111111111, 16'b1111111111111100, 16'b0000000000000000, 16'b0000000000000011, 16'b1111111111110100, 16'b0000000000010100, 16'b0000000000000100, 16'b0000000000011101, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000010101000, 16'b1111111111110001, 16'b1111111111111010, 16'b1111111111111111, 16'b1111111111100100, 16'b1111111111110101, 16'b0000000000101101}, 
{16'b0000000000001111, 16'b0000000000010010, 16'b0000000001010011, 16'b1111111111110101, 16'b0000000000011001, 16'b0000000001011001, 16'b0000000000000000, 16'b1111111111111000, 16'b0000000000011110, 16'b1111111111100010, 16'b1111111111111111, 16'b1111111111100001, 16'b0000000000000000, 16'b0000000001100100, 16'b1111111111111011, 16'b0000000000000000, 16'b0000000000111100, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111110101111, 16'b1111111111000001, 16'b1111111111110110, 16'b1111111111111111, 16'b1111111111011010, 16'b1111111111110110, 16'b1111111111101010, 16'b1111111111001101, 16'b1111111111001001, 16'b0000000000000111, 16'b0000000000011100, 16'b1111111110011010, 16'b0000000000000000}, 
{16'b1111111110110011, 16'b0000000000000000, 16'b1111111111111100, 16'b1111111111110011, 16'b1111111111111111, 16'b0000000000100010, 16'b1111111111101100, 16'b0000000001000101, 16'b1111111110100011, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111101000, 16'b0000000000010100, 16'b0000000000101110, 16'b1111111111111101, 16'b1111111110111111, 16'b1111111111110000, 16'b0000000000011100, 16'b0000000000010000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000010100, 16'b1111111111000010, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111011111}, 
{16'b1111111110101001, 16'b1111111111111110, 16'b1111111111111111, 16'b1111111111111011, 16'b1111111111111110, 16'b0000000000011011, 16'b0000000000000001, 16'b0000000000001000, 16'b0000000000001001, 16'b0000000000010000, 16'b0000000000010100, 16'b0000000000101001, 16'b0000000000000110, 16'b1111111111100111, 16'b0000000000000000, 16'b0000000001100001, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000011100, 16'b0000000000100100, 16'b0000000000000111, 16'b0000000000001010, 16'b1111111111111000, 16'b1111111111110111, 16'b0000000000000110, 16'b1111111111101110, 16'b1111111111011111, 16'b0000000000110101, 16'b1111111111111000, 16'b0000000000001000, 16'b1111111111001111}, 
{16'b0000000000000000, 16'b1111111111111111, 16'b0000000000001001, 16'b0000000000000000, 16'b0000000011101000, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000011100, 16'b1111111111101100, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000100001, 16'b0000000000000000, 16'b1111111111011010, 16'b1111111111111111, 16'b1111111111101110, 16'b0000000001010011, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000010001, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000001010}, 
{16'b1111111111111111, 16'b0000000000000111, 16'b1111111111111111, 16'b0000000000001100, 16'b1111111111110100, 16'b1111111111100001, 16'b1111111111110000, 16'b0000000001000111, 16'b0000000000000000, 16'b0000000000011000, 16'b1111111111111101, 16'b0000000000010000, 16'b1111111111110111, 16'b1111111111010111, 16'b1111111111001111, 16'b0000000000000011, 16'b1111111111111111, 16'b1111111111110111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000010011, 16'b0000000000001001, 16'b1111111111011111, 16'b0000000000011100, 16'b1111111111010101, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111010101, 16'b0000000000000000, 16'b0000000000001011, 16'b1111111111111000}, 
{16'b1111111111111101, 16'b1111111111100110, 16'b0000000000000000, 16'b1111111111110000, 16'b0000000000110111, 16'b1111111111111111, 16'b1111111111111010, 16'b0000000000011011, 16'b1111111110011011, 16'b0000000000000000, 16'b1111111111110110, 16'b1111111111111111, 16'b0000000001011001, 16'b0000000000111010, 16'b1111111111100110, 16'b1111111111111010, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111011101, 16'b1111111111100001, 16'b0000000000100001, 16'b0000000000000000, 16'b1111111111011100, 16'b0000000000000110, 16'b1111111111101011, 16'b1111111111110111, 16'b0000000000100010, 16'b0000000000000000, 16'b1111111111000000}, 
{16'b0000000010100010, 16'b0000000001010111, 16'b1111111111000000, 16'b0000000000000000, 16'b1111111110100111, 16'b0000000000000000, 16'b0000000000111001, 16'b0000000000000111, 16'b0000000000111001, 16'b1111111111111111, 16'b1111111111011000, 16'b1111111111101011, 16'b0000000000100100, 16'b0000000000000111, 16'b1111111111100110, 16'b0000000000100001, 16'b0000000010001001, 16'b1111111111011110, 16'b1111111110110100, 16'b0000000000000000, 16'b1111111111111000, 16'b1111111111010010, 16'b1111111111111100, 16'b1111111111111111, 16'b0000000000010110, 16'b1111111110100011, 16'b0000000000010110, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000011011, 16'b1111111111111000, 16'b0000000000001111}, 
{16'b1111111111101000, 16'b1111111111001110, 16'b1111111111110110, 16'b1111111111010101, 16'b1111111111111011, 16'b0000000000001100, 16'b0000000000000000, 16'b1111111111111101, 16'b0000000000001001, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111001000, 16'b0000000000011010, 16'b0000000000010100, 16'b1111111111100101, 16'b0000000001110001, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111110, 16'b0000000000000000, 16'b0000000001010000, 16'b1111111110000111, 16'b1111111111100100, 16'b1111111111110001, 16'b1111111111111011, 16'b0000000000110010, 16'b1111111111110010, 16'b0000000000000100, 16'b0000000001111011, 16'b1111111101111100, 16'b1111111110100010, 16'b0000000000000101}, 
{16'b0000000000000100, 16'b1111111111110000, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111101000111, 16'b1111111101100100, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111110111100, 16'b0000000000000110, 16'b0000000000000000, 16'b1111111111111000, 16'b0000000000000000, 16'b1111111111110001, 16'b1111111111110010, 16'b1111111111101110, 16'b1111111111011010, 16'b0000000001001000, 16'b0000000000000000, 16'b0000000000001011, 16'b1111111111111111, 16'b1111111111101101, 16'b0000000000000000, 16'b1111111111101001, 16'b0000000000111000, 16'b1111111101100000, 16'b0000000000111000, 16'b1111111111111111, 16'b1111111111111110, 16'b0000000000110011, 16'b1111111111111111, 16'b0000000000111100}, 
{16'b1111111111111111, 16'b0000000000000001, 16'b1111111111110100, 16'b0000000000010011, 16'b0000000000001110, 16'b1111111110101000, 16'b0000000000000000, 16'b0000000000010000, 16'b0000000010010100, 16'b1111111111111101, 16'b0000000000000000, 16'b0000000000001110, 16'b0000000001011011, 16'b1111111111110111, 16'b0000000000000011, 16'b0000000000011001, 16'b1111111111111111, 16'b0000000000000111, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111110111001, 16'b0000000000001001, 16'b0000000000010001, 16'b0000000000000101, 16'b1111111111111111, 16'b0000000000110111, 16'b0000000000000001, 16'b0000000000100000, 16'b1111111110010101, 16'b0000000000011010, 16'b0000000001100101, 16'b0000000000000001}, 
{16'b1111111110100110, 16'b0000000000110110, 16'b1111111110111101, 16'b0000000000011111, 16'b1111111111100101, 16'b0000000000000000, 16'b0000000001111111, 16'b1111111111000100, 16'b1111111110110101, 16'b0000000000101011, 16'b1111111111000110, 16'b1111111111111001, 16'b1111111111111111, 16'b0000000001011000, 16'b1111111111111111, 16'b1111111110110010, 16'b1111111111111111, 16'b0000000001110000, 16'b1111111110000111, 16'b1111111111111001, 16'b0000000001010001, 16'b1111111110100011, 16'b0000000000001101, 16'b1111111111111100, 16'b0000000001000101, 16'b1111111101111101, 16'b1111111110100011, 16'b1111111111001101, 16'b1111111111111111, 16'b0000000000011010, 16'b0000000000000110, 16'b0000000000101101}, 
{16'b1111111111101000, 16'b0000000000001101, 16'b1111111111111111, 16'b0000000000100110, 16'b1111111111110110, 16'b0000000000111010, 16'b0000000000000000, 16'b1111111111111101, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000010000101, 16'b0000000000000011, 16'b0000000000110000, 16'b0000000000000000, 16'b1111111111001001, 16'b1111111111101100, 16'b1111111111111111, 16'b1111111111111011, 16'b0000000000001010, 16'b1111111111111111, 16'b1111111111010000, 16'b1111111111111111, 16'b0000000001001011, 16'b0000000001001111, 16'b1111111111111111, 16'b1111111111111011, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111100111}, 
{16'b1111111111101011, 16'b0000000000000000, 16'b0000000001000101, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111100010, 16'b0000000000000000, 16'b1111111100100010, 16'b0000000000110111, 16'b0000000000000011, 16'b0000000000000110, 16'b1111111110100011, 16'b0000000000000000, 16'b1111111111011100, 16'b1111111111110111, 16'b0000000000000000, 16'b0000000000000101, 16'b0000000000000000, 16'b0000000000011100, 16'b0000000000000000, 16'b1111111111111101, 16'b0000000001010100, 16'b0000000001100000, 16'b1111111111000111, 16'b1111111111011011, 16'b0000000000111111, 16'b1111111110110001, 16'b0000000000000111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000101111}, 
{16'b1111111111100010, 16'b1111111111111111, 16'b1111111111000010, 16'b1111111111001100, 16'b1111111111111100, 16'b1111111111011101, 16'b0000000000000000, 16'b0000000000010111, 16'b1111111111000010, 16'b1111111111101010, 16'b1111111111110011, 16'b0000000000000000, 16'b0000000000000111, 16'b1111111111111101, 16'b1111111111110000, 16'b0000000000011000, 16'b0000000000111001, 16'b0000000000100001, 16'b1111111111011110, 16'b0000000000001100, 16'b1111111111111100, 16'b1111111111111000, 16'b0000000000000101, 16'b0000000000000100, 16'b1111111111101110, 16'b0000000000010110, 16'b1111111111101000, 16'b0000000000001111, 16'b1111111111111111, 16'b1111111110110100, 16'b1111111111111001, 16'b0000000000111001}, 
{16'b1111111111111001, 16'b1111111111101010, 16'b0000000000010011, 16'b0000000001000000, 16'b0000000000010101, 16'b0000000000010101, 16'b0000000000001011, 16'b1111111111001100, 16'b1111111111001011, 16'b0000000000010001, 16'b0000000000000011, 16'b0000000000001011, 16'b0000000000000101, 16'b0000000000000001, 16'b0000000000110100, 16'b0000000000000001, 16'b1111111111110010, 16'b0000000000011010, 16'b1111111111111000, 16'b1111111111110110, 16'b0000000000011100, 16'b1111111111100000, 16'b1111111111111001, 16'b0000000000100000, 16'b0000000000000101, 16'b1111111111100100, 16'b1111111111001101, 16'b1111111111111100, 16'b1111111110111000, 16'b0000000000001111, 16'b0000000000011010, 16'b0000000000000000}, 
{16'b1111111111111100, 16'b1111111111111010, 16'b1111111111111100, 16'b1111111111110111, 16'b1111111111011110, 16'b1111111111011100, 16'b0000000000010000, 16'b0000000000000010, 16'b1111111111010001, 16'b0000000000101010, 16'b1111111111111010, 16'b1111111111111111, 16'b1111111111100011, 16'b0000000000000001, 16'b0000000000000111, 16'b1111111111110010, 16'b1111111111111011, 16'b1111111111110101, 16'b1111111111101011, 16'b0000000000000000, 16'b1111111111011100, 16'b0000000000011010, 16'b1111111111001001, 16'b0000000000000001, 16'b0000000000001010, 16'b0000000000011111, 16'b0000000000000110, 16'b0000000000000001, 16'b0000000001001010, 16'b0000000000001101, 16'b0000000000000000, 16'b0000000000010101}, 
{16'b1111111111111011, 16'b0000000001000000, 16'b1111111111111111, 16'b1111111111110111, 16'b1111111111001001, 16'b1111111111101100, 16'b0000000001101001, 16'b1111111101001111, 16'b1111111110100110, 16'b1111111111001100, 16'b1111111111000111, 16'b1111111110111111, 16'b1111111111111111, 16'b0000000001111011, 16'b1111111111111001, 16'b0000000000000000, 16'b1111111111001001, 16'b0000000001110010, 16'b1111111110010110, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111110101001, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000001110, 16'b1111111111110001, 16'b1111111111011010, 16'b1111111111111111, 16'b0000000000101100, 16'b0000000000000000, 16'b1111111111101011, 16'b0000000000000000}, 
{16'b0000000001011110, 16'b1111111111100011, 16'b0000000000100001, 16'b1111111111110111, 16'b0000000000010011, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111101000, 16'b0000000000000000, 16'b0000000000010111, 16'b1111111111111111, 16'b1111111111110000, 16'b1111111111111111, 16'b0000000000111010, 16'b0000000000000100, 16'b0000000000001010, 16'b0000000000000110, 16'b1111111111111001, 16'b0000000000000101, 16'b0000000000000000, 16'b1111111111111101, 16'b1111111111111111, 16'b1111111110110001, 16'b1111111111111111, 16'b0000000000001110, 16'b1111111111100010, 16'b1111111111011101, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000010001110, 16'b1111111110110110, 16'b1111111111100010}, 
{16'b1111111111110100, 16'b1111111111100101, 16'b1111111111101111, 16'b0000000000001001, 16'b0000000000100011, 16'b1111111111011110, 16'b1111111111111111, 16'b1111111111000111, 16'b0000000000001111, 16'b0000000000100010, 16'b1111111111001001, 16'b1111111110111111, 16'b0000000000000110, 16'b1111111101010001, 16'b1111111111101100, 16'b1111111111100000, 16'b1111111111001101, 16'b1111111111111111, 16'b0000000000100010, 16'b0000000000000000, 16'b1111111111110100, 16'b1111111111110100, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111110000, 16'b1111111100111110, 16'b1111111101110001, 16'b1111111110111010, 16'b0000000000001110, 16'b0000000000110100, 16'b1111111111111111, 16'b0000000000111101}, 
{16'b1111111111101000, 16'b1111111111001001, 16'b0000000000101001, 16'b0000000000010011, 16'b0000000000001011, 16'b1111111111101000, 16'b1111111111110111, 16'b0000000000011001, 16'b0000000010001001, 16'b1111111111010100, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000011110, 16'b1111111111110001, 16'b1111111111111011, 16'b1111111111111011, 16'b1111111111100110, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000111010, 16'b1111111111011101, 16'b1111111111111111, 16'b0000000000100000, 16'b1111111111111101, 16'b0000000000000000, 16'b0000000010000110, 16'b0000000001010011, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111110010100, 16'b1111111111101110, 16'b1111111111111111}, 
{16'b0000000000000011, 16'b0000000000001100, 16'b1111111111111100, 16'b0000000000000000, 16'b0000000000111011, 16'b1111111110000100, 16'b0000000000000000, 16'b1111111111100111, 16'b0000000000101111, 16'b0000000000000000, 16'b1111111111111011, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000001, 16'b1111111111100100, 16'b0000000001000010, 16'b1111111111111110, 16'b1111111111111100, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111110, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000011, 16'b1111111110101110, 16'b0000000000001101, 16'b0000000000101110, 16'b1111111111111111, 16'b0000000000011000, 16'b1111111111111111, 16'b0000000000010011}, 
{16'b1111111111001100, 16'b0000000000000010, 16'b1111111110000100, 16'b0000000000000001, 16'b1111111111110011, 16'b1111111111110101, 16'b1111111111111111, 16'b1111111111101000, 16'b1111111111110110, 16'b1111111111101111, 16'b0000000000001100, 16'b0000000000000110, 16'b1111111111010010, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111101, 16'b0000000000010010, 16'b1111111111111010, 16'b1111111111111000, 16'b1111111111111000, 16'b1111111111111111, 16'b0000000001000101, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111101, 16'b0000000001010001, 16'b0000000000110000, 16'b0000000000001000, 16'b1111111111100111, 16'b1111111111111101, 16'b0000000000010000, 16'b0000000000001110}, 
{16'b0000000000001000, 16'b0000000000001010, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111110001000, 16'b0000000000001011, 16'b0000000000000110, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111010100, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111010110, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111110100100, 16'b0000000000000010, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000100001, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000001110100, 16'b0000000001010111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111000100, 16'b0000000000000000, 16'b1111111111111111}, 
{16'b0000000000010011, 16'b0000000000001101, 16'b0000000001000000, 16'b1111111111000000, 16'b0000000000100001, 16'b0000000000011110, 16'b0000000000000001, 16'b0000000000110001, 16'b0000000000000011, 16'b1111111111111100, 16'b0000000000001001, 16'b0000000000000001, 16'b1111111111111111, 16'b0000000000011110, 16'b1111111111111110, 16'b1111111111110101, 16'b0000000000000000, 16'b0000000000001000, 16'b1111111111110011, 16'b0000000000011001, 16'b0000000000001000, 16'b1111111101101011, 16'b1111111111100010, 16'b0000000000010111, 16'b1111111111111111, 16'b1111111101111110, 16'b1111111111011111, 16'b1111111111111010, 16'b1111111111111111, 16'b1111111111110001, 16'b0000000000000000, 16'b1111111111110101}, 
{16'b0000000000000000, 16'b1111111111111111, 16'b1111111111101000, 16'b1111111111010100, 16'b0000000000001010, 16'b0000000000000000, 16'b0000000000011000, 16'b1111111111111110, 16'b0000000000111111, 16'b1111111111111110, 16'b0000000000000000, 16'b1111111110101000, 16'b1111111111111111, 16'b0000000000100000, 16'b1111111111111111, 16'b1111111110111101, 16'b0000000000000000, 16'b1111111111111101, 16'b0000000001000011, 16'b1111111111111111, 16'b1111111110010000, 16'b1111111111111111, 16'b0000000001000010, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000100011, 16'b1111111111100111, 16'b0000000000010001, 16'b0000000000000000, 16'b1111111111001100, 16'b0000000000000000, 16'b0000000000000000}, 
{16'b1111111111001000, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111110, 16'b0000000001111110, 16'b1111111111100000, 16'b1111111111111110, 16'b1111111111111110, 16'b1111111111110100, 16'b1111111111110011, 16'b0000000000010000, 16'b0000000000100010, 16'b1111111111110110, 16'b0000000000111111, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111110110111, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111101011, 16'b0000000000000000, 16'b0000000000001001, 16'b0000000000000011, 16'b1111111111111101, 16'b1111111111110010, 16'b1111111111001100, 16'b1111111110110100, 16'b0000000000000000, 16'b1111111111100011, 16'b0000000000001010, 16'b1111111111111111, 16'b0000000000010011}, 
{16'b1111111110010110, 16'b1111111111010111, 16'b1111111111011000, 16'b0000000000000000, 16'b0000000010010010, 16'b1111111111000111, 16'b0000000000000000, 16'b1111111111110010, 16'b1111111110010111, 16'b0000000000100011, 16'b1111111111111111, 16'b0000000010010001, 16'b0000000000000000, 16'b1111111111110011, 16'b1111111111111111, 16'b0000000000001000, 16'b1111111111111011, 16'b0000000000000000, 16'b1111111111110100, 16'b0000000001111110, 16'b0000000000001001, 16'b1111111111110101, 16'b0000000000011100, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111100111, 16'b1111111111110100, 16'b1111111110001000, 16'b1111111111011011, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111110000}, 
{16'b0000000000111001, 16'b1111111100110011, 16'b1111111101000110, 16'b1111111111010100, 16'b0000000010101011, 16'b1111111111111111, 16'b1111111110100111, 16'b0000000001000011, 16'b0000000000001111, 16'b0000000000000000, 16'b0000000000110101, 16'b1111111110111010, 16'b0000000000000000, 16'b0000000000000001, 16'b1111111111110111, 16'b0000000000000100, 16'b1111111111100101, 16'b1111111100010100, 16'b0000000000101010, 16'b0000000001011000, 16'b0000000001000011, 16'b0000000000000000, 16'b0000000000000111, 16'b1111111110011000, 16'b1111111101011110, 16'b1111111111111110, 16'b1111111110110011, 16'b1111111110001010, 16'b1111111111001110, 16'b1111111100011111, 16'b0000000001101011, 16'b0000000001101101}, 
{16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000001000010, 16'b1111111111010000, 16'b0000000000000100, 16'b0000000000010010, 16'b1111111110100110, 16'b0000000000001001, 16'b1111111111111110, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000111101, 16'b0000000000001101, 16'b0000000000000101, 16'b0000000000001111, 16'b0000000001010101, 16'b1111111111001000, 16'b0000000000000000, 16'b1111111111010101, 16'b1111111111111111, 16'b0000000001010000, 16'b0000000000000010, 16'b1111111111111111, 16'b1111111101110000, 16'b1111111111111101, 16'b1111111111011000, 16'b1111111111110000, 16'b0000000000000000, 16'b0000000000100010, 16'b0000000000011010}, 
{16'b1111111111110100, 16'b0000000000100010, 16'b1111111110110010, 16'b0000000000000101, 16'b0000000000110001, 16'b1111111111110101, 16'b1111111111111110, 16'b0000000000101001, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111101111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111110111, 16'b1111111111100000, 16'b1111111111101111, 16'b1111111111110001, 16'b1111111111101111, 16'b1111111111100011, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111110100, 16'b1111111111101110, 16'b0000000001100101, 16'b0000000000000000, 16'b1111111110100011, 16'b1111111111111101, 16'b0000000000011111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000001000000, 16'b1111111111111111}, 
{16'b1111111111111111, 16'b0000000000000001, 16'b1111111111111111, 16'b1111111111011000, 16'b1111111100100011, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111110, 16'b1111111101100110, 16'b0000000000010100, 16'b1111111111100110, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111110100001, 16'b1111111111110100, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000010, 16'b0000000000001001, 16'b0000000001011000, 16'b1111111111100001, 16'b1111111110110011, 16'b0000000000000000, 16'b1111111110111101, 16'b1111111111100110, 16'b1111111111000100, 16'b1111111111111110, 16'b1111111111111100, 16'b1111111111111011, 16'b1111111110000111, 16'b1111111111110111, 16'b0000000000111110}, 
{16'b0000000000011100, 16'b0000000000111000, 16'b1111111111111111, 16'b0000000000101000, 16'b1111111111001010, 16'b1111111111100000, 16'b0000000000011000, 16'b0000000000010001, 16'b1111111111110011, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111110101101, 16'b1111111111111111, 16'b0000000000100100, 16'b1111111111100010, 16'b0000000000001000, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000110101, 16'b1111111110101100, 16'b0000000001000111, 16'b0000000000001100, 16'b0000000000000000, 16'b0000000000110110, 16'b0000000000000000, 16'b1111111111110110, 16'b1111111110011110, 16'b1111111111100011, 16'b1111111111010100, 16'b0000000000101101}, 
{16'b0000000000000000, 16'b0000000000000001, 16'b1111111110100010, 16'b1111111111111111, 16'b0000000000110100, 16'b1111111111011011, 16'b1111111111111100, 16'b1111111111111111, 16'b0000000000000101, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111001011, 16'b0000000000011000, 16'b0000000000000001, 16'b0000000000000000, 16'b0000000000001001, 16'b1111111111111111, 16'b1111111111011001, 16'b0000000000000100, 16'b0000000000000000, 16'b1111111111110111, 16'b1111111111111010, 16'b0000000001001011, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111110110101, 16'b1111111110101100, 16'b0000000000111101, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000111, 16'b0000000001001000}, 
{16'b1111111110101000, 16'b1111111111111111, 16'b1111111111001001, 16'b0000000000000001, 16'b1111111110100101, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111101111, 16'b1111111101110111, 16'b1111111111111001, 16'b0000000000000000, 16'b1111111111111101, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111101, 16'b1111111111110011, 16'b1111111111011010, 16'b1111111111100111, 16'b0000000000010000, 16'b1111111111111111, 16'b1111111111111001, 16'b0000000000000000, 16'b0000000001010110, 16'b1111111111111111, 16'b0000000000100110, 16'b0000000000010111, 16'b1111111111011100, 16'b0000000000110110, 16'b1111111111110100, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000010010101}, 
{16'b1111111110101111, 16'b0000000000000111, 16'b0000000000001100, 16'b1111111111111000, 16'b0000000000111110, 16'b1111111110110010, 16'b1111111111111110, 16'b0000000001000011, 16'b0000000000101000, 16'b0000000000000010, 16'b1111111111111111, 16'b1111111111101110, 16'b1111111111101001, 16'b1111111111101111, 16'b1111111111110011, 16'b0000000000010111, 16'b1111111111111111, 16'b0000000000000010, 16'b0000000000100100, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000011, 16'b0000000001000000, 16'b0000000000001011, 16'b0000000000000001, 16'b1111111111100100, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111100, 16'b1111111111111100, 16'b1111111111111111, 16'b0000000000010001}, 
{16'b1111111111111111, 16'b0000000000000000, 16'b1111111111001001, 16'b1111111111101100, 16'b0000000001001000, 16'b1111111111111111, 16'b1111111111101100, 16'b0000000000111110, 16'b1111111111110010, 16'b0000000001001010, 16'b0000000000010101, 16'b1111111111100001, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111100, 16'b0000000000000101, 16'b1111111111101100, 16'b1111111110111100, 16'b0000000001000111, 16'b0000000000100111, 16'b0000000010100010, 16'b0000000000110011, 16'b0000000000111111, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000001110, 16'b0000000000010100, 16'b1111111110010100, 16'b1111111111111111, 16'b1111111111111110, 16'b1111111111111110}, 
{16'b0000000000000000, 16'b1111111111101001, 16'b1111111111100101, 16'b0000000000000000, 16'b1111111111000001, 16'b0000000000000000, 16'b0000000000110001, 16'b0000000000011011, 16'b0000000000001101, 16'b1111111111100110, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111110101, 16'b0000000000110011, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111110110010, 16'b0000000000000000, 16'b1111111111001110, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111110, 16'b0000000000000011, 16'b0000000000000100, 16'b0000000000000111, 16'b0000000000100011, 16'b1111111111101111, 16'b1111111111111110, 16'b1111111110001101, 16'b0000000000010100}, 
{16'b0000000001110001, 16'b1111111111111101, 16'b0000000000010000, 16'b1111111111100101, 16'b1111111111101010, 16'b0000000000001000, 16'b0000000000101001, 16'b0000000000000000, 16'b0000000010000110, 16'b0000000000000000, 16'b1111111111111010, 16'b0000000000000100, 16'b0000000000011000, 16'b1111111111111111, 16'b0000000000001101, 16'b0000000000011010, 16'b1111111111111110, 16'b1111111110001110, 16'b1111111111110001, 16'b1111111111111111, 16'b0000000000011101, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000011100, 16'b0000000000000100, 16'b1111111110111100, 16'b1111111111100101, 16'b0000000000100001, 16'b1111111111111000, 16'b0000000001000010, 16'b1111111111111111, 16'b1111111111010010}, 
{16'b0000000000000011, 16'b0000000000011010, 16'b1111111111111111, 16'b1111111111110110, 16'b1111111110100101, 16'b1111111111111111, 16'b0000000000001011, 16'b1111111111110100, 16'b0000000000101010, 16'b1111111111110111, 16'b1111111111111111, 16'b1111111111110111, 16'b1111111111111111, 16'b1111111111110110, 16'b0000000000000000, 16'b0000000001010000, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000001000, 16'b0000000000100000, 16'b0000000000000000, 16'b0000000000000001, 16'b0000000000001000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000101, 16'b0000000000000000, 16'b0000000000011000}, 
{16'b1111111110110000, 16'b0000000000100001, 16'b0000000000000100, 16'b1111111111100101, 16'b1111111110011001, 16'b1111111111111011, 16'b0000000000010001, 16'b1111111110011010, 16'b0000000010000010, 16'b0000000000010010, 16'b0000000000000100, 16'b0000000000011000, 16'b0000000000001011, 16'b0000000000000000, 16'b0000000001101000, 16'b1111111111101010, 16'b0000000000000001, 16'b0000000000000000, 16'b1111111111111110, 16'b0000000000000000, 16'b1111111110010001, 16'b0000000000000100, 16'b0000000000100111, 16'b0000000000001001, 16'b0000000000001001, 16'b1111111101010111, 16'b1111111110101000, 16'b1111111111000010, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000001010011, 16'b1111111111001011}, 
{16'b1111111111111100, 16'b1111111111001110, 16'b1111111111100101, 16'b1111111110010111, 16'b1111111110111101, 16'b0000000001010110, 16'b0000000001001111, 16'b1111111111010100, 16'b0000000000001010, 16'b1111111111110110, 16'b1111111111100111, 16'b1111111110111111, 16'b0000000000011010, 16'b1111111110110111, 16'b0000000000110000, 16'b1111111111111111, 16'b0000000001010101, 16'b1111111111111111, 16'b1111111111111110, 16'b1111111111011101, 16'b1111111111110101, 16'b1111111111101111, 16'b1111111110111011, 16'b0000000000010101, 16'b1111111111111111, 16'b1111111111111110, 16'b1111111111000101, 16'b0000000001010000, 16'b0000000001000111, 16'b1111111111101000, 16'b1111111101011110, 16'b0000000000100100}, 
{16'b0000000000000000, 16'b1111111111111001, 16'b1111111111111111, 16'b1111111111100111, 16'b0000000000000111, 16'b0000000000000010, 16'b0000000000010001, 16'b0000000000000001, 16'b0000000000011110, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000011000, 16'b0000000000000000, 16'b0000000000000011, 16'b1111111111011110, 16'b1111111111100100, 16'b0000000000000000, 16'b0000000000101110, 16'b0000000000001110, 16'b0000000000100000, 16'b1111111111111011, 16'b1111111111010111, 16'b1111111111111111, 16'b0000000000010011, 16'b1111111111111111, 16'b0000000000001000, 16'b1111111111111110, 16'b0000000000010001, 16'b0000000000000000, 16'b0000000000010101, 16'b1111111110011110, 16'b1111111111111111}, 
{16'b0000000001001111, 16'b1111111111111101, 16'b0000000000100110, 16'b1111111110110001, 16'b1111111111001110, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000111, 16'b0000000000000000, 16'b1111111111011111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111011110, 16'b0000000000100100, 16'b1111111111111111, 16'b1111111111111000, 16'b0000000000000000, 16'b0000000000011110, 16'b1111111111001100, 16'b0000000000011101, 16'b0000000000100011, 16'b0000000000100001, 16'b1111111111111111, 16'b0000000010001101, 16'b1111111111011000, 16'b0000000001011101, 16'b1111111111110010, 16'b1111111110100011, 16'b1111111111010011, 16'b0000000000100011}, 
{16'b1111111101110100, 16'b1111111111111001, 16'b1111111111011000, 16'b1111111111111111, 16'b0000000001000010, 16'b1111111111010010, 16'b1111111111110000, 16'b0000000000111100, 16'b0000000000011000, 16'b1111111111000011, 16'b0000000000000000, 16'b1111111111111000, 16'b1111111111111101, 16'b0000000000100011, 16'b1111111111000001, 16'b1111111111111101, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111011, 16'b0000000000000000, 16'b1111111111001111, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111110101011, 16'b0000000000010001, 16'b0000000010011110, 16'b0000000001011000, 16'b1111111111110110, 16'b1111111111010110, 16'b1111111110001101, 16'b0000000000000000, 16'b1111111111110011}, 
{16'b0000000000000101, 16'b0000000000110110, 16'b0000000000000101, 16'b1111111111011001, 16'b0000000000000001, 16'b1111111111111001, 16'b0000000000000000, 16'b0000000000110101, 16'b0000000000110111, 16'b1111111111011101, 16'b0000000000100011, 16'b0000000000000110, 16'b1111111111111111, 16'b1111111111111100, 16'b1111111111010111, 16'b0000000001000000, 16'b1111111111110101, 16'b1111111110101101, 16'b0000000000011101, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000011101, 16'b1111111111101100, 16'b1111111111111110, 16'b1111111111110010, 16'b0000000000010110, 16'b1111111111011100, 16'b0000000000100010, 16'b1111111110100010, 16'b0000000000010100, 16'b1111111111111111, 16'b0000000000101000}, 
{16'b1111111111110101, 16'b0000000000000000, 16'b0000000000010110, 16'b0000000000000000, 16'b1111111111110000, 16'b1111111111111111, 16'b0000000000011010, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000001, 16'b0000000000000000, 16'b0000000000000101, 16'b1111111111100100, 16'b0000000000000010, 16'b0000000000011100, 16'b0000000000001011, 16'b0000000000011011, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000100000, 16'b0000000000111111, 16'b1111111111100110, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000010, 16'b1111111110001001, 16'b1111111111111111, 16'b1111111111101101, 16'b1111111111111111, 16'b0000000010010000, 16'b0000000000000000, 16'b1111111111001011}, 
{16'b1111111111111001, 16'b1111111111100001, 16'b1111111111111101, 16'b0000000000000001, 16'b0000000000010111, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111010, 16'b0000000000010010, 16'b1111111111111101, 16'b0000000000000000, 16'b0000000000001000, 16'b0000000001001011, 16'b1111111111100101, 16'b0000000000000011, 16'b1111111100100110, 16'b1111111111111101, 16'b1111111111110000, 16'b0000000000000010, 16'b1111111111110011, 16'b0000000000010111, 16'b1111111111000110, 16'b0000000000011101, 16'b0000000000011010, 16'b1111111111111100, 16'b1111111101001001, 16'b1111111111000101, 16'b1111111111111010, 16'b1111111111111011, 16'b0000000001100011, 16'b1111111111111110, 16'b0000000000100111}, 
{16'b0000000000001100, 16'b0000000000000000, 16'b0000000000101100, 16'b1111111111100010, 16'b1111111111101110, 16'b0000000000111100, 16'b1111111111010111, 16'b0000000000001110, 16'b1111111110110000, 16'b0000000000000010, 16'b0000000000000100, 16'b1111111111101010, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111001111, 16'b0000000001101110, 16'b1111111111000000, 16'b1111111111111100, 16'b0000000000011110, 16'b1111111111111111, 16'b0000000000010001, 16'b1111111110000101, 16'b0000000001010000, 16'b1111111111111111, 16'b1111111111100000, 16'b0000000001111100, 16'b0000000000100101, 16'b1111111111010111, 16'b1111111111011101, 16'b1111111101110110, 16'b1111111111111101, 16'b0000000000000100}, 
{16'b1111111111111111, 16'b0000000000000001, 16'b1111111111110111, 16'b1111111110111011, 16'b1111111111111111, 16'b1111111110011011, 16'b0000000000000000, 16'b0000000001001101, 16'b0000000000111110, 16'b0000000000000100, 16'b0000000000000000, 16'b1111111111100011, 16'b0000000001010101, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000001101111, 16'b0000000000000000, 16'b1111111111110101, 16'b1111111111110010, 16'b1111111110101101, 16'b0000000000100001, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000001000, 16'b1111111111101101, 16'b1111111110001010, 16'b0000000001000110, 16'b1111111110001110, 16'b0000000000001101, 16'b1111111111101011, 16'b0000000000000000}, 
{16'b0000000000001111, 16'b0000000000101111, 16'b0000000000000010, 16'b1111111111111111, 16'b1111111110001010, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000111110, 16'b0000000001000110, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000101011, 16'b1111111111100101, 16'b1111111110010001, 16'b1111111111110111, 16'b1111111111100110, 16'b1111111111100111, 16'b1111111111101110, 16'b1111111111111111, 16'b1111111111101111, 16'b1111111111111010, 16'b1111111111111101, 16'b0000000000100100, 16'b1111111111111111, 16'b0000000001110110}
};

localparam logic signed [15:0] bias [32] = '{
16'b0000000101111001,  // 1.474280834197998
16'b0000000010110001,  // 0.6914801001548767
16'b0000000101110000,  // 1.4406442642211914
16'b0000000101101000,  // 1.408045768737793
16'b0000000011111100,  // 0.9864811301231384
16'b0000000011011101,  // 0.8636202812194824
16'b1111111101100010,  // -0.6153604388237
16'b0000000001111011,  // 0.4839226007461548
16'b0000000001111100,  // 0.4862793982028961
16'b0000000001011111,  // 0.37162142992019653
16'b0000000001110101,  // 0.45989668369293213
16'b0000000101001100,  // 1.2998151779174805
16'b1111111011111011,  // -1.016528844833374
16'b1111111110100101,  // -0.35249894857406616
16'b0000000001110010,  // 0.44582197070121765
16'b1111111111100011,  // -0.1119980737566948
16'b1111111111101110,  // -0.06717441976070404
16'b0000000000000001,  // 0.00487547367811203
16'b0000000000110001,  // 0.1946917623281479
16'b1111111100111000,  // -0.7796769738197327
16'b0000000010111010,  // 0.7287401556968689
16'b0000000110110111,  // 1.714877724647522
16'b1111111001100111,  // -1.5971007347106934
16'b0000000000010010,  // 0.07393483817577362
16'b0000000001010010,  // 0.3225609362125397
16'b0000000011011000,  // 0.8453295230865479
16'b0000000011100110,  // 0.898597240447998
16'b0000000001000001,  // 0.2548799514770508
16'b0000000011111001,  // 0.9735668301582336
16'b0000000100100000,  // 1.1261906623840332
16'b0000000001110010,  // 0.44768181443214417
16'b1111110110100001   // -2.3676068782806396
};
endpackage