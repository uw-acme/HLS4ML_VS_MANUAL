package softmax_invert_16_10;
localparam logic signed invert_table = {
16'h1FFFF,
16'h01000,
16'h00800,
16'h00555,
16'h00400,
16'h00333,
16'h002AB,
16'h00249,
16'h00200,
16'h001C7,
16'h0019A,
16'h00174,
16'h00155,
16'h0013B,
16'h00125,
16'h00111,
16'h00100,
16'h000F1,
16'h000E4,
16'h000D8,
16'h000CD,
16'h000C3,
16'h000BA,
16'h000B2,
16'h000AB,
16'h000A4,
16'h0009E,
16'h00098,
16'h00092,
16'h0008D,
16'h00089,
16'h00084,
16'h00080,
16'h0007C,
16'h00078,
16'h00075,
16'h00072,
16'h0006F,
16'h0006C,
16'h00069,
16'h00066,
16'h00064,
16'h00062,
16'h0005F,
16'h0005D,
16'h0005B,
16'h00059,
16'h00057,
16'h00055,
16'h00054,
16'h00052,
16'h00050,
16'h0004F,
16'h0004D,
16'h0004C,
16'h0004A,
16'h00049,
16'h00048,
16'h00047,
16'h00045,
16'h00044,
16'h00043,
16'h00042,
16'h00041,
16'h00040,
16'h0003F,
16'h0003E,
16'h0003D,
16'h0003C,
16'h0003B,
16'h0003B,
16'h0003A,
16'h00039,
16'h00038,
16'h00037,
16'h00037,
16'h00036,
16'h00035,
16'h00035,
16'h00034,
16'h00033,
16'h00033,
16'h00032,
16'h00031,
16'h00031,
16'h00030,
16'h00030,
16'h0002F,
16'h0002F,
16'h0002E,
16'h0002E,
16'h0002D,
16'h0002D,
16'h0002C,
16'h0002C,
16'h0002B,
16'h0002B,
16'h0002A,
16'h0002A,
16'h00029,
16'h00029,
16'h00029,
16'h00028,
16'h00028,
16'h00027,
16'h00027,
16'h00027,
16'h00026,
16'h00026,
16'h00026,
16'h00025,
16'h00025,
16'h00025,
16'h00024,
16'h00024,
16'h00024,
16'h00023,
16'h00023,
16'h00023,
16'h00022,
16'h00022,
16'h00022,
16'h00022,
16'h00021,
16'h00021,
16'h00021,
16'h00021,
16'h00020,
16'h00020,
16'h00020,
16'h00020,
16'h0001F,
16'h0001F,
16'h0001F,
16'h0001F,
16'h0001E,
16'h0001E,
16'h0001E,
16'h0001E,
16'h0001D,
16'h0001D,
16'h0001D,
16'h0001D,
16'h0001D,
16'h0001C,
16'h0001C,
16'h0001C,
16'h0001C,
16'h0001C,
16'h0001B,
16'h0001B,
16'h0001B,
16'h0001B,
16'h0001B,
16'h0001B,
16'h0001A,
16'h0001A,
16'h0001A,
16'h0001A,
16'h0001A,
16'h0001A,
16'h00019,
16'h00019,
16'h00019,
16'h00019,
16'h00019,
16'h00019,
16'h00019,
16'h00018,
16'h00018,
16'h00018,
16'h00018,
16'h00018,
16'h00018,
16'h00018,
16'h00017,
16'h00017,
16'h00017,
16'h00017,
16'h00017,
16'h00017,
16'h00017,
16'h00017,
16'h00016,
16'h00016,
16'h00016,
16'h00016,
16'h00016,
16'h00016,
16'h00016,
16'h00016,
16'h00015,
16'h00015,
16'h00015,
16'h00015,
16'h00015,
16'h00015,
16'h00015,
16'h00015,
16'h00015,
16'h00014,
16'h00014,
16'h00014,
16'h00014,
16'h00014,
16'h00014,
16'h00014,
16'h00014,
16'h00014,
16'h00014,
16'h00014,
16'h00013,
16'h00013,
16'h00013,
16'h00013,
16'h00013,
16'h00013,
16'h00013,
16'h00013,
16'h00013,
16'h00013,
16'h00013,
16'h00012,
16'h00012,
16'h00012,
16'h00012,
16'h00012,
16'h00012,
16'h00012,
16'h00012,
16'h00012,
16'h00012,
16'h00012,
16'h00012,
16'h00012,
16'h00011,
16'h00011,
16'h00011,
16'h00011,
16'h00011,
16'h00011,
16'h00011,
16'h00011,
16'h00011,
16'h00011,
16'h00011,
16'h00011,
16'h00011,
16'h00011,
16'h00010,
16'h00010,
16'h00010,
16'h00010,
16'h00010,
16'h00010,
16'h00010,
16'h00010,
16'h00010,
16'h00010,
16'h00010,
16'h00010,
16'h00010,
16'h00010,
16'h00010,
16'h00010,
16'h0000F,
16'h0000F,
16'h0000F,
16'h0000F,
16'h0000F,
16'h0000F,
16'h0000F,
16'h0000F,
16'h0000F,
16'h0000F,
16'h0000F,
16'h0000F,
16'h0000F,
16'h0000F,
16'h0000F,
16'h0000F,
16'h0000F,
16'h0000F,
16'h0000E,
16'h0000E,
16'h0000E,
16'h0000E,
16'h0000E,
16'h0000E,
16'h0000E,
16'h0000E,
16'h0000E,
16'h0000E,
16'h0000E,
16'h0000E,
16'h0000E,
16'h0000E,
16'h0000E,
16'h0000E,
16'h0000E,
16'h0000E,
16'h0000E,
16'h0000E,
16'h0000E,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000D,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000C,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000B,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h0000A,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00009,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h00008,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF8,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF7,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF6,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF5,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF4,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF3,
16'h3FFF2,
16'h3FFF2,
16'h3FFF2,
16'h3FFF2,
16'h3FFF2,
16'h3FFF2,
16'h3FFF2,
16'h3FFF2,
16'h3FFF2,
16'h3FFF2,
16'h3FFF2,
16'h3FFF2,
16'h3FFF2,
16'h3FFF2,
16'h3FFF2,
16'h3FFF2,
16'h3FFF2,
16'h3FFF2,
16'h3FFF2,
16'h3FFF2,
16'h3FFF2,
16'h3FFF1,
16'h3FFF1,
16'h3FFF1,
16'h3FFF1,
16'h3FFF1,
16'h3FFF1,
16'h3FFF1,
16'h3FFF1,
16'h3FFF1,
16'h3FFF1,
16'h3FFF1,
16'h3FFF1,
16'h3FFF1,
16'h3FFF1,
16'h3FFF1,
16'h3FFF1,
16'h3FFF1,
16'h3FFF1,
16'h3FFF0,
16'h3FFF0,
16'h3FFF0,
16'h3FFF0,
16'h3FFF0,
16'h3FFF0,
16'h3FFF0,
16'h3FFF0,
16'h3FFF0,
16'h3FFF0,
16'h3FFF0,
16'h3FFF0,
16'h3FFF0,
16'h3FFF0,
16'h3FFF0,
16'h3FFF0,
16'h3FFEF,
16'h3FFEF,
16'h3FFEF,
16'h3FFEF,
16'h3FFEF,
16'h3FFEF,
16'h3FFEF,
16'h3FFEF,
16'h3FFEF,
16'h3FFEF,
16'h3FFEF,
16'h3FFEF,
16'h3FFEF,
16'h3FFEF,
16'h3FFEE,
16'h3FFEE,
16'h3FFEE,
16'h3FFEE,
16'h3FFEE,
16'h3FFEE,
16'h3FFEE,
16'h3FFEE,
16'h3FFEE,
16'h3FFEE,
16'h3FFEE,
16'h3FFEE,
16'h3FFEE,
16'h3FFED,
16'h3FFED,
16'h3FFED,
16'h3FFED,
16'h3FFED,
16'h3FFED,
16'h3FFED,
16'h3FFED,
16'h3FFED,
16'h3FFED,
16'h3FFED,
16'h3FFEC,
16'h3FFEC,
16'h3FFEC,
16'h3FFEC,
16'h3FFEC,
16'h3FFEC,
16'h3FFEC,
16'h3FFEC,
16'h3FFEC,
16'h3FFEC,
16'h3FFEC,
16'h3FFEB,
16'h3FFEB,
16'h3FFEB,
16'h3FFEB,
16'h3FFEB,
16'h3FFEB,
16'h3FFEB,
16'h3FFEB,
16'h3FFEB,
16'h3FFEA,
16'h3FFEA,
16'h3FFEA,
16'h3FFEA,
16'h3FFEA,
16'h3FFEA,
16'h3FFEA,
16'h3FFEA,
16'h3FFE9,
16'h3FFE9,
16'h3FFE9,
16'h3FFE9,
16'h3FFE9,
16'h3FFE9,
16'h3FFE9,
16'h3FFE9,
16'h3FFE8,
16'h3FFE8,
16'h3FFE8,
16'h3FFE8,
16'h3FFE8,
16'h3FFE8,
16'h3FFE8,
16'h3FFE7,
16'h3FFE7,
16'h3FFE7,
16'h3FFE7,
16'h3FFE7,
16'h3FFE7,
16'h3FFE7,
16'h3FFE6,
16'h3FFE6,
16'h3FFE6,
16'h3FFE6,
16'h3FFE6,
16'h3FFE6,
16'h3FFE5,
16'h3FFE5,
16'h3FFE5,
16'h3FFE5,
16'h3FFE5,
16'h3FFE5,
16'h3FFE4,
16'h3FFE4,
16'h3FFE4,
16'h3FFE4,
16'h3FFE4,
16'h3FFE3,
16'h3FFE3,
16'h3FFE3,
16'h3FFE3,
16'h3FFE3,
16'h3FFE2,
16'h3FFE2,
16'h3FFE2,
16'h3FFE2,
16'h3FFE1,
16'h3FFE1,
16'h3FFE1,
16'h3FFE1,
16'h3FFE0,
16'h3FFE0,
16'h3FFE0,
16'h3FFE0,
16'h3FFDF,
16'h3FFDF,
16'h3FFDF,
16'h3FFDF,
16'h3FFDE,
16'h3FFDE,
16'h3FFDE,
16'h3FFDE,
16'h3FFDD,
16'h3FFDD,
16'h3FFDD,
16'h3FFDC,
16'h3FFDC,
16'h3FFDC,
16'h3FFDB,
16'h3FFDB,
16'h3FFDB,
16'h3FFDA,
16'h3FFDA,
16'h3FFDA,
16'h3FFD9,
16'h3FFD9,
16'h3FFD9,
16'h3FFD8,
16'h3FFD8,
16'h3FFD7,
16'h3FFD7,
16'h3FFD7,
16'h3FFD6,
16'h3FFD6,
16'h3FFD5,
16'h3FFD5,
16'h3FFD4,
16'h3FFD4,
16'h3FFD3,
16'h3FFD3,
16'h3FFD2,
16'h3FFD2,
16'h3FFD1,
16'h3FFD1,
16'h3FFD0,
16'h3FFD0,
16'h3FFCF,
16'h3FFCF,
16'h3FFCE,
16'h3FFCD,
16'h3FFCD,
16'h3FFCC,
16'h3FFCB,
16'h3FFCB,
16'h3FFCA,
16'h3FFC9,
16'h3FFC9,
16'h3FFC8,
16'h3FFC7,
16'h3FFC6,
16'h3FFC5,
16'h3FFC5,
16'h3FFC4,
16'h3FFC3,
16'h3FFC2,
16'h3FFC1,
16'h3FFC0,
16'h3FFBF,
16'h3FFBE,
16'h3FFBD,
16'h3FFBC,
16'h3FFBB,
16'h3FFB9,
16'h3FFB8,
16'h3FFB7,
16'h3FFB6,
16'h3FFB4,
16'h3FFB3,
16'h3FFB1,
16'h3FFB0,
16'h3FFAE,
16'h3FFAC,
16'h3FFAB,
16'h3FFA9,
16'h3FFA7,
16'h3FFA5,
16'h3FFA3,
16'h3FFA1,
16'h3FF9E,
16'h3FF9C,
16'h3FF9A,
16'h3FF97,
16'h3FF94,
16'h3FF91,
16'h3FF8E,
16'h3FF8B,
16'h3FF88,
16'h3FF84,
16'h3FF80,
16'h3FF7C,
16'h3FF77,
16'h3FF73,
16'h3FF6E,
16'h3FF68,
16'h3FF62,
16'h3FF5C,
16'h3FF55,
16'h3FF4E,
16'h3FF46,
16'h3FF3D,
16'h3FF33,
16'h3FF28,
16'h3FF1C,
16'h3FF0F,
16'h3FF00,
16'h3FEEF,
16'h3FEDB,
16'h3FEC5,
16'h3FEAB,
16'h3FE8C,
16'h3FE66,
16'h3FE39,
16'h3FE00,
16'h3FDB7,
16'h3FD55,
16'h3FCCD,
16'h3FC00,
16'h3FAAB,
16'h3F800,
16'h3F000,
};
endpackage