// Width: 19
// NFRAC: 10
package dense_4_19_10;

localparam logic signed [18:0] weights [32][5] = '{ 
{19'b1111111111111110011, 19'b0000000000101000011, 19'b1111111111011001110, 19'b0000000000001000011, 19'b1111111111110010011}, 
{19'b1111111110111000100, 19'b1111111111111000111, 19'b0000000000111010111, 19'b1111111111111110011, 19'b0000000000000010001}, 
{19'b0000000000101111100, 19'b0000000000011011000, 19'b1111111111111100011, 19'b1111111111001100000, 19'b1111111111100101000}, 
{19'b1111111111001111111, 19'b1111111111010000010, 19'b1111111111110001101, 19'b0000000000100111011, 19'b0000000000011110000}, 
{19'b0000000000001111101, 19'b0000000000010000011, 19'b0000000000010100000, 19'b1111111111111101101, 19'b1111111101111110010}, 
{19'b0000000000101001110, 19'b1111111111001101100, 19'b0000000000010111001, 19'b1111111111101011010, 19'b1111111111101010001}, 
{19'b1111111111001100101, 19'b0000000000000100100, 19'b1111111111111111111, 19'b0000000000010110010, 19'b0000000000001000110}, 
{19'b1111111111111111110, 19'b0000000000100100011, 19'b1111111111001101110, 19'b0000000000010100110, 19'b0000000000010001011}, 
{19'b0000000000010100111, 19'b1111111111101010010, 19'b0000000000000000001, 19'b1111111111000100111, 19'b1111111111100000001}, 
{19'b1111111111111111111, 19'b1111111111011101111, 19'b0000000000010110110, 19'b0000000000110111000, 19'b0000000000000000000}, 
{19'b1111111111101111010, 19'b1111111111101101011, 19'b0000000000000000000, 19'b0000000001001010011, 19'b1111111111011101101}, 
{19'b0000000000010101101, 19'b0000000000011101010, 19'b1111111111010100011, 19'b1111111111111100011, 19'b0000000000001111100}, 
{19'b0000000000000000000, 19'b0000000000010101011, 19'b0000000000000001001, 19'b1111111111100101011, 19'b1111111110110000010}, 
{19'b0000000000010110101, 19'b0000000000001000001, 19'b0000000000110101101, 19'b1111111111110111000, 19'b1111111111001001001}, 
{19'b0000000000001011100, 19'b1111111111111001110, 19'b1111111111010001110, 19'b1111111111111011110, 19'b0000000001000100101}, 
{19'b1111111111000011010, 19'b1111111111100000101, 19'b1111111111100011100, 19'b0000000000110011000, 19'b0000000000000100000}, 
{19'b0000000000101100010, 19'b1111111111101010000, 19'b1111111111101110101, 19'b1111111111100011000, 19'b1111111111111000010}, 
{19'b0000000000011000111, 19'b1111111111111010110, 19'b1111111111001011001, 19'b1111111111111100000, 19'b0000000000001001000}, 
{19'b0000000000100001000, 19'b0000000000000101010, 19'b1111111111100100000, 19'b0000000000000000000, 19'b1111111111001111111}, 
{19'b0000000000011101100, 19'b1111111111110100111, 19'b1111111111100100110, 19'b0000000000011010100, 19'b0000000000001100001}, 
{19'b0000000000001000101, 19'b1111111111111100000, 19'b0000000000100110000, 19'b1111111111001000110, 19'b1111111111111101010}, 
{19'b0000000000000000000, 19'b0000000000001111000, 19'b0000000000111110010, 19'b1111111110111101101, 19'b1111111110110000111}, 
{19'b1111111111110011011, 19'b0000000000001110000, 19'b0000000000010110101, 19'b1111111111010010010, 19'b0000000001000010110}, 
{19'b1111111111111111111, 19'b0000000000010101000, 19'b0000000000100100001, 19'b0000000000000100110, 19'b1111111110110110110}, 
{19'b1111111111101010010, 19'b0000000000101110101, 19'b1111111111100011011, 19'b0000000000000000101, 19'b0000000000110001101}, 
{19'b0000000000000011010, 19'b0000000000100010000, 19'b0000000000000011110, 19'b1111111110100000010, 19'b0000000001000110001}, 
{19'b1111111111000101001, 19'b1111111111100000110, 19'b0000000000011011011, 19'b0000000000011111010, 19'b0000000000011001110}, 
{19'b0000000000000000100, 19'b0000000000011110110, 19'b1111111111111011010, 19'b1111111111101100101, 19'b0000000000000100000}, 
{19'b1111111111110010101, 19'b0000000000011111100, 19'b1111111110111111100, 19'b0000000000010001110, 19'b1111111111101011101}, 
{19'b1111111111111101101, 19'b0000000000010010000, 19'b1111111111101010011, 19'b1111111111001100101, 19'b0000000001001011111}, 
{19'b0000000000111001011, 19'b0000000000001000111, 19'b0000000000101001100, 19'b1111111110110100100, 19'b1111111111010111101}, 
{19'b1111111111111000011, 19'b1111111111001110100, 19'b0000000000101110110, 19'b0000000000001001000, 19'b0000000000010000010}
};

localparam logic signed [18:0] bias [5] = '{
19'b1111111111111000000,  // -0.06223141402006149
19'b1111111111110111111,  // -0.06270556896924973
19'b1111111111110111000,  // -0.07014333456754684
19'b0000000000001010100,  // 0.0820775106549263
19'b0000000000011011100   // 0.2155742198228836
};
endpackage