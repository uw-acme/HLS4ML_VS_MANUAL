// Width: 22
// NFRAC: 11
package dense_2_22_11;

localparam logic signed [21:0] weights [64][32] = '{ 
{22'b0000000000001000100110, 22'b0000000000000000010000, 22'b1111111111111001111011, 22'b1111111111111111010100, 22'b0000000000001000010110, 22'b0000000000000000000000, 22'b1111111111111011011000, 22'b1111111111111111111111, 22'b1111111111110111001111, 22'b0000000000000010100011, 22'b0000000000000000000000, 22'b1111111111111111110100, 22'b1111111111111111111111, 22'b1111111111111001100110, 22'b1111111111111110011000, 22'b1111111111110111100111, 22'b0000000000000000000000, 22'b1111111111111111100101, 22'b1111111111111001111001, 22'b1111111111111010111011, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b1111111111111111101111, 22'b1111111111111111111010, 22'b0000000000000000000000, 22'b0000000000000011001101, 22'b0000000000001100010110, 22'b0000000000000101100110, 22'b1111111111111111111111, 22'b0000000000000001100111, 22'b1111111111110010111001, 22'b0000000000000000000000}, 
{22'b1111111111111100110010, 22'b1111111111111011000010, 22'b1111111111111011100100, 22'b1111111111111110001110, 22'b1111111111111111110100, 22'b0000000000000001011000, 22'b1111111111111000110110, 22'b0000000000000000001010, 22'b0000000000000000001001, 22'b1111111111111101111111, 22'b0000000000000100111111, 22'b1111111111111110100111, 22'b1111111111111110000111, 22'b1111111111111001000011, 22'b0000000000000000001111, 22'b1111111111111110011101, 22'b0000000000000000011001, 22'b1111111111111001110001, 22'b0000000000000101011111, 22'b0000000000000111010110, 22'b1111111111111110111111, 22'b1111111111111111110100, 22'b1111111111111111111111, 22'b0000000000000000110000, 22'b1111111111111101101110, 22'b0000000000001000110011, 22'b0000000000000111111011, 22'b0000000000000000010001, 22'b0000000000000000111010, 22'b1111111111110000011011, 22'b0000000000000000001111, 22'b0000000000000000000000}, 
{22'b0000000000000010010100, 22'b1111111111111100010101, 22'b1111111111111011110110, 22'b1111111111111110101010, 22'b1111111111111101100001, 22'b1111111111111101010001, 22'b1111111111111010000101, 22'b0000000000000000001001, 22'b1111111111111011101011, 22'b0000000000000000010010, 22'b0000000000000000000100, 22'b1111111111111101011010, 22'b0000000000000010111001, 22'b1111111111111101111011, 22'b1111111111111111111101, 22'b1111111111111110110100, 22'b0000000000000000001010, 22'b0000000000000011000011, 22'b0000000000000001111000, 22'b0000000000000111010110, 22'b0000000000000001010100, 22'b1111111111111101010011, 22'b0000000000000000000000, 22'b0000000000000001000111, 22'b1111111111111111011010, 22'b0000000000000110101100, 22'b0000000000000100110001, 22'b0000000000000011000110, 22'b1111111111111111111111, 22'b1111111111111011001000, 22'b1111111111111111100100, 22'b0000000000000011001011}, 
{22'b0000000000000100011010, 22'b0000000000000000100111, 22'b0000000000000001101100, 22'b1111111111111111101100, 22'b1111111111101111101101, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b0000000000000111001111, 22'b0000000000000111110000, 22'b1111111111111111100100, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b0000000000000000001010, 22'b1111111111111111011010, 22'b0000000000000110110111, 22'b0000000000000000000000, 22'b1111111111111111001101, 22'b1111111111111111111111, 22'b1111111111111010010111, 22'b1111111111111110000010, 22'b0000000000000001100101, 22'b1111111111111101111110, 22'b1111111111111111111111, 22'b0000000000000000000111, 22'b1111111111111110011000, 22'b0000000000000010010101, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b1111111111111001000111, 22'b0000000000001001111011}, 
{22'b1111111111101010001010, 22'b1111111111111111001101, 22'b1111111111111111110111, 22'b0000000000000000001010, 22'b1111111111111111001010, 22'b0000000000000000001101, 22'b1111111111111110011011, 22'b1111111111111011001101, 22'b0000000000000001101111, 22'b1111111111111111010110, 22'b1111111111111111100100, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b0000000000000110101110, 22'b0000000000000000000000, 22'b0000000000001010100001, 22'b1111111111111111111111, 22'b0000000000000110111110, 22'b1111111111110011001100, 22'b0000000000000000000000, 22'b1111111111111100011011, 22'b0000000000000101011001, 22'b0000000000001000010000, 22'b0000000000000000000000, 22'b0000000000000001011100, 22'b0000000000000101001101, 22'b0000000000000111101000, 22'b0000000000000000100011, 22'b1111111111111111110110, 22'b1111111111111111111111, 22'b1111111111111111100011, 22'b0000000000000111001111}, 
{22'b0000000000000001110110, 22'b1111111111111111111111, 22'b0000000000000100110001, 22'b1111111111101011001111, 22'b1111111111010011111011, 22'b1111111111110100110010, 22'b0000000000001011010101, 22'b1111111111101100000101, 22'b1111111111111111111111, 22'b1111111111101010010100, 22'b1111111111101111111101, 22'b1111111111110101000101, 22'b0000000000001011010011, 22'b1111111111111111111111, 22'b1111111111111111100001, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b1111111111111011110001, 22'b1111111111111111111111, 22'b1111111111110000010110, 22'b0000000000000000000000, 22'b0000000000000101111100, 22'b1111111111111111111111, 22'b0000000000000000101101, 22'b0000000000001000100100, 22'b0000000000000001101000, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b0000000000000110100101, 22'b1111111111111110111010, 22'b0000000000000110011010}, 
{22'b1111111111111110110110, 22'b1111111111111010111101, 22'b1111111111111000010001, 22'b1111111111111110011111, 22'b1111111111110110110001, 22'b0000000000000010000111, 22'b1111111111111010001111, 22'b1111111111111011011101, 22'b1111111111110010101110, 22'b0000000000000001100011, 22'b1111111111111111110101, 22'b1111111111111010111010, 22'b0000000000000011110011, 22'b1111111111111111101011, 22'b1111111111111110101011, 22'b1111111111101110010010, 22'b1111111111111111111111, 22'b0000000000000010101100, 22'b0000000000000110001000, 22'b1111111111111010110011, 22'b1111111111111011001100, 22'b1111111111111101111111, 22'b1111111111111111111101, 22'b0000000000000000111000, 22'b1111111111111110100010, 22'b1111111111101011010000, 22'b1111111111110111100001, 22'b1111111111111110100011, 22'b0000000000000000001011, 22'b1111111111111111010100, 22'b0000000000000000111110, 22'b1111111111111111111110}, 
{22'b1111111111111011000101, 22'b1111111111111101000110, 22'b1111111111111101011101, 22'b1111111111111000011010, 22'b1111111111111100010010, 22'b1111111111111111111111, 22'b0000000000000011010101, 22'b1111111111111101011110, 22'b0000000000000110011010, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b0000000000000111000000, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b1111111111111101101111, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b1111111111111111111110, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b0000000000000001011010, 22'b1111111111111010001111, 22'b0000000000000000011100, 22'b1111111111111111111111, 22'b1111111111111101101100, 22'b1111111111111111111110, 22'b0000000000000000000000, 22'b1111111111111111111111}, 
{22'b1111111111110000101110, 22'b1111111111111110001011, 22'b1111111111110011110101, 22'b0000000000000011111010, 22'b0000000000001111100101, 22'b1111111111111111111111, 22'b1111111111111111000100, 22'b0000000000000111101001, 22'b1111111111110001111101, 22'b1111111111111110100000, 22'b0000000000000000000000, 22'b1111111111111001100011, 22'b1111111111111111111111, 22'b0000000000000010011011, 22'b1111111111111001111001, 22'b0000000000011000001000, 22'b1111111111111111101110, 22'b0000000000000001011111, 22'b0000000000000110101001, 22'b0000000000000111110101, 22'b0000000000000000000000, 22'b1111111111110101010000, 22'b0000000000000000000000, 22'b0000000000001101001010, 22'b1111111111111010001100, 22'b0000000000010110010100, 22'b1111111111111011001110, 22'b1111111111111001011110, 22'b1111111111110000111001, 22'b1111111111110001001001, 22'b0000000000000000000000, 22'b0000000000000001101101}, 
{22'b0000000000000000000000, 22'b1111111111111111100000, 22'b1111111111111101101000, 22'b0000000000000000000000, 22'b0000000000001001110111, 22'b1111111111111111010110, 22'b1111111111111101111101, 22'b0000000000000010111100, 22'b0000000000000011001111, 22'b0000000000000000000111, 22'b1111111111111111101110, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b1111111111111100010111, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b1111111111111111110101, 22'b0000000000000000000100, 22'b0000000000000010101101, 22'b0000000000000000100111, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b0000000000000000001110, 22'b0000000000000001001110, 22'b1111111111111011110001, 22'b0000000000000010001011, 22'b0000000000000111111101, 22'b1111111111111111111111, 22'b0000000000000000001100, 22'b0000000000000001100101, 22'b0000000000000010001110}, 
{22'b0000000000000011000101, 22'b0000000000000000000000, 22'b1111111111111100101100, 22'b1111111111110111111110, 22'b1111111111100110100101, 22'b0000000000000100010000, 22'b0000000000000000000000, 22'b1111111111100101100001, 22'b0000000000000001001010, 22'b1111111111111111111111, 22'b0000000000000000000111, 22'b1111111111111111111100, 22'b0000000000000000010101, 22'b0000000000000000000000, 22'b1111111111111111011001, 22'b1111111111110011110010, 22'b1111111111111111111111, 22'b0000000000000111000010, 22'b0000000000000100000010, 22'b0000000000000110000111, 22'b1111111111110001111011, 22'b1111111111110100100111, 22'b0000000000000011110101, 22'b1111111111111110111000, 22'b1111111111111110100001, 22'b0000000000001011011110, 22'b1111111111111100111010, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b0000000000000110110000, 22'b1111111111111111111111, 22'b0000000000000000001100}, 
{22'b1111111111111001101011, 22'b1111111111110000001110, 22'b0000000000000000000000, 22'b1111111111111111111011, 22'b0000000000001010101000, 22'b1111111111110111011000, 22'b1111111111111000111010, 22'b0000000000000011101101, 22'b1111111111111111111110, 22'b0000000000000100110000, 22'b0000000000000010010111, 22'b1111111111111101100101, 22'b0000000000000000000000, 22'b0000000000000000011100, 22'b1111111111111111010100, 22'b1111111111110111111001, 22'b0000000000000101100111, 22'b0000000000000000111010, 22'b0000000000001001100000, 22'b0000000000000010110001, 22'b0000000000000000000000, 22'b1111111111111110110010, 22'b0000000000000100000010, 22'b1111111111111101001111, 22'b1111111111110110001001, 22'b1111111111111111110010, 22'b0000000000000101111010, 22'b1111111111111111111111, 22'b0000000000000000010001, 22'b1111111111111100111110, 22'b0000000000000100011001, 22'b0000000000001000110101}, 
{22'b0000000000000000011111, 22'b0000000000000000000000, 22'b0000000000000111000001, 22'b0000000000000000010001, 22'b1111111111111110101100, 22'b0000000000000101110001, 22'b0000000000000010111100, 22'b1111111111111111111111, 22'b0000000000000000000001, 22'b1111111111111011100000, 22'b1111111111111110010000, 22'b1111111111111010101001, 22'b1111111111111111111111, 22'b0000000000000001100111, 22'b1111111111111101110010, 22'b0000000000011010111110, 22'b0000000000000000000000, 22'b1111111111111100111111, 22'b1111111111111001111101, 22'b1111111111111111100100, 22'b0000000000000110010110, 22'b0000000000000100000110, 22'b0000000000000000000000, 22'b1111111111111111111010, 22'b0000000000000111000001, 22'b0000000000001000100101, 22'b0000000000001111110110, 22'b0000000000000000010101, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b1111111111111111100111, 22'b1111111111111101101101}, 
{22'b1111111111111011000000, 22'b0000000000000001100011, 22'b0000000000000001010000, 22'b1111111111111000000101, 22'b1111111111110111011000, 22'b0000000000001111000000, 22'b0000000000000001100100, 22'b0000000000000000000000, 22'b1111111111111010110110, 22'b1111111111111101001011, 22'b0000000000000100001001, 22'b0000000000000010010001, 22'b0000000000000000000001, 22'b1111111111111101011111, 22'b0000000000001001001001, 22'b1111111111111111111111, 22'b1111111111111111100100, 22'b0000000000000000000000, 22'b0000000000000000011010, 22'b1111111111111110100000, 22'b0000000000000010100000, 22'b0000000000000000100000, 22'b0000000000000011101001, 22'b1111111111111111111111, 22'b0000000000000000000110, 22'b0000000000010101000011, 22'b1111111111111110001100, 22'b1111111111111111010000, 22'b1111111111111111111111, 22'b1111111111111100100000, 22'b1111111111111110101101, 22'b0000000000000101101000}, 
{22'b0000000000000001111000, 22'b0000000000000010010111, 22'b0000000000001010011100, 22'b1111111111111110101110, 22'b0000000000000011001110, 22'b0000000000001011001110, 22'b0000000000000000000001, 22'b1111111111111111000011, 22'b0000000000000011110001, 22'b1111111111111100010110, 22'b1111111111111111111111, 22'b1111111111111100001011, 22'b0000000000000000000000, 22'b0000000000001100100101, 22'b1111111111111111011011, 22'b0000000000000000000011, 22'b0000000000000111100011, 22'b0000000000000000000001, 22'b0000000000000000000110, 22'b1111111111110101111111, 22'b1111111111111000001001, 22'b1111111111111110110110, 22'b1111111111111111111111, 22'b1111111111111011010101, 22'b1111111111111110110110, 22'b1111111111111101010111, 22'b1111111111111001101101, 22'b1111111111111001001100, 22'b0000000000000000111101, 22'b0000000000000011100100, 22'b1111111111110011010010, 22'b0000000000000000000110}, 
{22'b1111111111110110011100, 22'b0000000000000000000000, 22'b1111111111111111100001, 22'b1111111111111110011010, 22'b1111111111111111111111, 22'b0000000000000100010001, 22'b1111111111111101100001, 22'b0000000000001000101011, 22'b1111111111110100011000, 22'b1111111111111111111110, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b1111111111111111111000, 22'b1111111111111101000110, 22'b0000000000000010100010, 22'b0000000000000101110111, 22'b1111111111111111101100, 22'b1111111111110111111101, 22'b1111111111111110000111, 22'b0000000000000011100101, 22'b0000000000000010000001, 22'b0000000000000000000000, 22'b0000000000000000000110, 22'b0000000000000010100111, 22'b1111111111111000010101, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b0000000000000000000110, 22'b0000000000000000000001, 22'b1111111111111011111110}, 
{22'b1111111111110101001111, 22'b1111111111111111110100, 22'b1111111111111111111001, 22'b1111111111111111011100, 22'b1111111111111111110110, 22'b0000000000000011011000, 22'b0000000000000000001101, 22'b0000000000000001000110, 22'b0000000000000001001110, 22'b0000000000000010000000, 22'b0000000000000010100001, 22'b0000000000000101001010, 22'b0000000000000000110110, 22'b1111111111111100111001, 22'b0000000000000000000001, 22'b0000000000001100001101, 22'b0000000000000000000000, 22'b0000000000000000000010, 22'b1111111111111111111010, 22'b0000000000000011100001, 22'b0000000000000100100011, 22'b0000000000000000111111, 22'b0000000000000001010100, 22'b1111111111111111000011, 22'b1111111111111110111110, 22'b0000000000000000110110, 22'b1111111111111101110110, 22'b1111111111111011111100, 22'b0000000000000110101101, 22'b1111111111111111000001, 22'b0000000000000001000000, 22'b1111111111111001111111}, 
{22'b0000000000000000000000, 22'b1111111111111111111111, 22'b0000000000000001001101, 22'b0000000000000000000000, 22'b0000000000011101000000, 22'b1111111111111111111110, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b0000000000000011100000, 22'b1111111111111101100110, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b0000000000000000000010, 22'b0000000000000100001000, 22'b0000000000000000000000, 22'b1111111111111011010110, 22'b1111111111111111111111, 22'b1111111111111101110110, 22'b0000000000001010011110, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b0000000000000010001011, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b0000000000000001010100}, 
{22'b1111111111111111111001, 22'b0000000000000000111011, 22'b1111111111111111111110, 22'b0000000000000001100010, 22'b1111111111111110100101, 22'b1111111111111100001011, 22'b1111111111111110000000, 22'b0000000000001000111000, 22'b0000000000000000000000, 22'b0000000000000011000110, 22'b1111111111111111101001, 22'b0000000000000010000100, 22'b1111111111111110111100, 22'b1111111111111010111101, 22'b1111111111111001111001, 22'b0000000000000000011010, 22'b1111111111111111111111, 22'b1111111111111110111000, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b1111111111111111111110, 22'b0000000000000010011011, 22'b0000000000000001001001, 22'b1111111111111011111110, 22'b0000000000000011100100, 22'b1111111111111010101111, 22'b0000000000000000000100, 22'b0000000000000000000000, 22'b1111111111111010101000, 22'b0000000000000000000000, 22'b0000000000000001011101, 22'b1111111111111111000000}, 
{22'b1111111111111111101000, 22'b1111111111111100110101, 22'b0000000000000000000000, 22'b1111111111111110000101, 22'b0000000000000110111010, 22'b1111111111111111111111, 22'b1111111111111111010101, 22'b0000000000000011011010, 22'b1111111111110011011111, 22'b0000000000000000000000, 22'b1111111111111110110001, 22'b1111111111111111111011, 22'b0000000000001011001111, 22'b0000000000000111010101, 22'b1111111111111100110100, 22'b1111111111111111010101, 22'b1111111111111111111111, 22'b0000000000000000000001, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b1111111111111011101001, 22'b1111111111111100001100, 22'b0000000000000100001100, 22'b0000000000000000000000, 22'b1111111111111011100111, 22'b0000000000000000110010, 22'b1111111111111101011011, 22'b1111111111111110111011, 22'b0000000000000100010110, 22'b0000000000000000000001, 22'b1111111111111000000101}, 
{22'b0000000000010100010011, 22'b0000000000001010111100, 22'b1111111111111000000001, 22'b0000000000000000000110, 22'b1111111111110100111011, 22'b0000000000000000000000, 22'b0000000000000111001000, 22'b0000000000000000111111, 22'b0000000000000111001010, 22'b1111111111111111111111, 22'b1111111111111011000010, 22'b1111111111111101011111, 22'b0000000000000100100010, 22'b0000000000000000111000, 22'b1111111111111100110110, 22'b0000000000000100001101, 22'b0000000000010001001000, 22'b1111111111111011110101, 22'b1111111111110110100001, 22'b0000000000000000000000, 22'b1111111111111111000101, 22'b1111111111111010010110, 22'b1111111111111111100111, 22'b1111111111111111111100, 22'b0000000000000010110000, 22'b1111111111110100011101, 22'b0000000000000010110110, 22'b1111111111111111111101, 22'b0000000000000000000000, 22'b0000000000000011011111, 22'b1111111111111111000100, 22'b0000000000000001111010}, 
{22'b1111111111111101000010, 22'b1111111111111001110110, 22'b1111111111111110110101, 22'b1111111111111010101001, 22'b1111111111111111011100, 22'b0000000000000001100100, 22'b0000000000000000000000, 22'b1111111111111111101000, 22'b0000000000000001001101, 22'b1111111111111111111000, 22'b0000000000000000000000, 22'b1111111111111001000011, 22'b0000000000000011010000, 22'b0000000000000010100100, 22'b1111111111111100101110, 22'b0000000000001110001100, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b1111111111111111110111, 22'b0000000000000000000000, 22'b0000000000001010000111, 22'b1111111111110000111100, 22'b1111111111111100100010, 22'b1111111111111110001101, 22'b1111111111111111011001, 22'b0000000000000110010011, 22'b1111111111111110010100, 22'b0000000000000000100100, 22'b0000000000001111011111, 22'b1111111111101111100110, 22'b1111111111110100010000, 22'b0000000000000000101101}, 
{22'b0000000000000000100010, 22'b1111111111111110000111, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b1111111111101000111111, 22'b1111111111101100100110, 22'b0000000000000000000011, 22'b1111111111111111111111, 22'b1111111111110111100001, 22'b0000000000000000110010, 22'b0000000000000000000000, 22'b1111111111111111000111, 22'b0000000000000000000000, 22'b1111111111111110001000, 22'b1111111111111110010100, 22'b1111111111111101110010, 22'b1111111111111011010010, 22'b0000000000001001000010, 22'b0000000000000000000000, 22'b0000000000000001011110, 22'b1111111111111111111111, 22'b1111111111111101101111, 22'b0000000000000000000000, 22'b1111111111111101001110, 22'b0000000000000111000001, 22'b1111111111101100000101, 22'b0000000000000111000010, 22'b1111111111111111111111, 22'b1111111111111111110110, 22'b0000000000000110011001, 22'b1111111111111111111111, 22'b0000000000000111100011}, 
{22'b1111111111111111111111, 22'b0000000000000000001010, 22'b1111111111111110100111, 22'b0000000000000010011001, 22'b0000000000000001110001, 22'b1111111111110101000011, 22'b0000000000000000000000, 22'b0000000000000010000011, 22'b0000000000010010100011, 22'b1111111111111111101101, 22'b0000000000000000000000, 22'b0000000000000001110011, 22'b0000000000001011011111, 22'b1111111111111110111110, 22'b0000000000000000011100, 22'b0000000000000011001110, 22'b1111111111111111111111, 22'b0000000000000000111000, 22'b1111111111111111111111, 22'b0000000000000000000001, 22'b1111111111110111001111, 22'b0000000000000001001110, 22'b0000000000000010001111, 22'b0000000000000000101110, 22'b1111111111111111111111, 22'b0000000000000110111111, 22'b0000000000000000001001, 22'b0000000000000100000010, 22'b1111111111110010101000, 22'b0000000000000011010010, 22'b0000000000001100101010, 22'b0000000000000000001011}, 
{22'b1111111111110100110001, 22'b0000000000000110110000, 22'b1111111111110111101010, 22'b0000000000000011111011, 22'b1111111111111100101000, 22'b0000000000000000000000, 22'b0000000000001111111011, 22'b1111111111111000100011, 22'b1111111111110110101011, 22'b0000000000000101011110, 22'b1111111111111000110111, 22'b1111111111111111001111, 22'b1111111111111111111110, 22'b0000000000001011000000, 22'b1111111111111111111100, 22'b1111111111110110010110, 22'b1111111111111111111111, 22'b0000000000001110000110, 22'b1111111111110000111011, 22'b1111111111111111001110, 22'b0000000000001010001000, 22'b1111111111110100011001, 22'b0000000000000001101100, 22'b1111111111111111100001, 22'b0000000000001000101011, 22'b1111111111101111101110, 22'b1111111111110100011001, 22'b1111111111111001101110, 22'b1111111111111111111111, 22'b0000000000000011010100, 22'b0000000000000000110011, 22'b0000000000000101101101}, 
{22'b1111111111111101000110, 22'b0000000000000001101010, 22'b1111111111111111111111, 22'b0000000000000100110010, 22'b1111111111111110110010, 22'b0000000000000111010000, 22'b0000000000000000000100, 22'b1111111111111111101001, 22'b1111111111111111111011, 22'b0000000000000000000010, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b1111111111111111111100, 22'b0000000000010000101001, 22'b0000000000000000011001, 22'b0000000000000110000010, 22'b0000000000000000000000, 22'b1111111111111001001110, 22'b1111111111111101100011, 22'b1111111111111111111111, 22'b1111111111111111011110, 22'b0000000000000001010110, 22'b1111111111111111111111, 22'b1111111111111010000100, 22'b1111111111111111111111, 22'b0000000000001001011101, 22'b0000000000001001111011, 22'b1111111111111111111111, 22'b1111111111111111011110, 22'b0000000000000000000000, 22'b1111111111111111111110, 22'b1111111111111100111010}, 
{22'b1111111111111101011010, 22'b0000000000000000000000, 22'b0000000000001000101111, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b1111111111111100010111, 22'b0000000000000000000000, 22'b1111111111100100010111, 22'b0000000000000110111001, 22'b0000000000000000011100, 22'b0000000000000000110110, 22'b1111111111110100011111, 22'b0000000000000000000110, 22'b1111111111111011100110, 22'b1111111111111110111100, 22'b0000000000000000000000, 22'b0000000000000000101000, 22'b0000000000000000000000, 22'b0000000000000011100110, 22'b0000000000000000000000, 22'b1111111111111111101101, 22'b0000000000001010100010, 22'b0000000000001100000011, 22'b1111111111111000111011, 22'b1111111111111011011101, 22'b0000000000000111111111, 22'b1111111111110110001110, 22'b0000000000000000111100, 22'b1111111111111111111110, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b0000000000000101111001}, 
{22'b1111111111111100010111, 22'b1111111111111111111110, 22'b1111111111111000010110, 22'b1111111111111001100010, 22'b1111111111111111100011, 22'b1111111111111011101011, 22'b0000000000000000000000, 22'b0000000000000010111010, 22'b1111111111111000010101, 22'b1111111111111101010101, 22'b1111111111111110011010, 22'b0000000000000000000000, 22'b0000000000000000111001, 22'b1111111111111111101011, 22'b1111111111111110000011, 22'b0000000000000011000011, 22'b0000000000000111001000, 22'b0000000000000100001100, 22'b1111111111111011110100, 22'b0000000000000001100011, 22'b1111111111111111100111, 22'b1111111111111111000101, 22'b0000000000000000101110, 22'b0000000000000000100000, 22'b1111111111111101110001, 22'b0000000000000010110110, 22'b1111111111111101000110, 22'b0000000000000001111010, 22'b1111111111111111111111, 22'b1111111111110110100011, 22'b1111111111111111001010, 22'b0000000000000111001100}, 
{22'b1111111111111111001000, 22'b1111111111111101010110, 22'b0000000000000010011101, 22'b0000000000001000000110, 22'b0000000000000010101101, 22'b0000000000000010101000, 22'b0000000000000001011111, 22'b1111111111111001100011, 22'b1111111111111001011011, 22'b0000000000000010001100, 22'b0000000000000000011000, 22'b0000000000000001011000, 22'b0000000000000000101101, 22'b0000000000000000001011, 22'b0000000000000110100100, 22'b0000000000000000001111, 22'b1111111111111110010001, 22'b0000000000000011010011, 22'b1111111111111111000011, 22'b1111111111111110110110, 22'b0000000000000011100001, 22'b1111111111111100000010, 22'b1111111111111111001001, 22'b0000000000000100000100, 22'b0000000000000000101101, 22'b1111111111111100100101, 22'b1111111111111001101010, 22'b1111111111111111100111, 22'b1111111111110111000100, 22'b0000000000000001111011, 22'b0000000000000011010000, 22'b0000000000000000000010}, 
{22'b1111111111111111100100, 22'b1111111111111111010111, 22'b1111111111111111100111, 22'b1111111111111110111001, 22'b1111111111111011110010, 22'b1111111111111011100000, 22'b0000000000000010000001, 22'b0000000000000000010000, 22'b1111111111111010001010, 22'b0000000000000101010110, 22'b1111111111111111010101, 22'b1111111111111111111110, 22'b1111111111111100011110, 22'b0000000000000000001010, 22'b0000000000000000111100, 22'b1111111111111110010100, 22'b1111111111111111011111, 22'b1111111111111110101010, 22'b1111111111111101011011, 22'b0000000000000000000000, 22'b1111111111111011100000, 22'b0000000000000011010000, 22'b1111111111111001001110, 22'b0000000000000000001010, 22'b0000000000000001010101, 22'b0000000000000011111101, 22'b0000000000000000110110, 22'b0000000000000000001100, 22'b0000000000001001010110, 22'b0000000000000001101001, 22'b0000000000000000000000, 22'b0000000000000010101011}, 
{22'b1111111111111111011000, 22'b0000000000001000000101, 22'b1111111111111111111111, 22'b1111111111111110111100, 22'b1111111111111001001010, 22'b1111111111111101100110, 22'b0000000000001101001010, 22'b1111111111101001111100, 22'b1111111111110100110100, 22'b1111111111111001100111, 22'b1111111111111000111110, 22'b1111111111110111111000, 22'b1111111111111111111110, 22'b0000000000001111011111, 22'b1111111111111111001010, 22'b0000000000000000000000, 22'b1111111111111001001111, 22'b0000000000001110010000, 22'b1111111111110010110010, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b1111111111110101001111, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b0000000000000001110011, 22'b1111111111111110001010, 22'b1111111111111011010001, 22'b1111111111111111111111, 22'b0000000000000101100101, 22'b0000000000000000000110, 22'b1111111111111101011011, 22'b0000000000000000000001}, 
{22'b0000000000001011110001, 22'b1111111111111100011010, 22'b0000000000000100001110, 22'b1111111111111110111101, 22'b0000000000000010011100, 22'b1111111111111111111000, 22'b1111111111111111111010, 22'b1111111111111101000001, 22'b0000000000000000000000, 22'b0000000000000010111100, 22'b1111111111111111111111, 22'b1111111111111110000111, 22'b1111111111111111111111, 22'b0000000000000111010100, 22'b0000000000000000100111, 22'b0000000000000001010010, 22'b0000000000000000110001, 22'b1111111111111111001110, 22'b0000000000000000101001, 22'b0000000000000000000000, 22'b1111111111111111101101, 22'b1111111111111111111111, 22'b1111111111110110001110, 22'b1111111111111111111111, 22'b0000000000000001110110, 22'b1111111111111100010001, 22'b1111111111111011101011, 22'b1111111111111111111111, 22'b1111111111111111111110, 22'b0000000000010001110110, 22'b1111111111110110110110, 22'b1111111111111100010010}, 
{22'b1111111111111110100101, 22'b1111111111111100101100, 22'b1111111111111101111011, 22'b0000000000000001001010, 22'b0000000000000100011101, 22'b1111111111111011110110, 22'b1111111111111111111101, 22'b1111111111111000111101, 22'b0000000000000001111100, 22'b0000000000000100010110, 22'b1111111111111001001010, 22'b1111111111110111111010, 22'b0000000000000000110000, 22'b1111111111101010001000, 22'b1111111111111101100101, 22'b1111111111111100000011, 22'b1111111111111001101010, 22'b1111111111111111111111, 22'b0000000000000100010010, 22'b0000000000000000000000, 22'b1111111111111110100010, 22'b1111111111111110100100, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b1111111111111110000111, 22'b1111111111100111110111, 22'b1111111111101110001110, 22'b1111111111110111010001, 22'b0000000000000001110010, 22'b0000000000000110100110, 22'b1111111111111111111111, 22'b0000000000000111101100}, 
{22'b1111111111111101000011, 22'b1111111111111001001000, 22'b0000000000000101001111, 22'b0000000000000010011000, 22'b0000000000000001011000, 22'b1111111111111101000011, 22'b1111111111111110111101, 22'b0000000000000011001001, 22'b0000000000010001001111, 22'b1111111111111010100001, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b0000000000000011110000, 22'b1111111111111110001111, 22'b1111111111111111011011, 22'b1111111111111111011101, 22'b1111111111111100110011, 22'b1111111111111111111110, 22'b0000000000000000000000, 22'b0000000000000111010000, 22'b1111111111111011101111, 22'b1111111111111111111001, 22'b0000000000000100000111, 22'b1111111111111111101011, 22'b0000000000000000000000, 22'b0000000000010000110101, 22'b0000000000001010011000, 22'b0000000000000000000110, 22'b0000000000000000000000, 22'b1111111111110010100010, 22'b1111111111111101110100, 22'b1111111111111111111111}, 
{22'b0000000000000000011110, 22'b0000000000000001100010, 22'b1111111111111111100011, 22'b0000000000000000000000, 22'b0000000000000111011001, 22'b1111111111110000100010, 22'b0000000000000000000000, 22'b1111111111111100111101, 22'b0000000000000101111101, 22'b0000000000000000000000, 22'b1111111111111111011010, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b0000000000000000001011, 22'b1111111111111100100011, 22'b0000000000001000010011, 22'b1111111111111111110100, 22'b1111111111111111100000, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b1111111111111111110000, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b0000000000000000011010, 22'b1111111111110101110110, 22'b0000000000000001101001, 22'b0000000000000101110111, 22'b1111111111111111111001, 22'b0000000000000011000001, 22'b1111111111111111111111, 22'b0000000000000010011001}, 
{22'b1111111111111001100011, 22'b0000000000000000010010, 22'b1111111111110000100100, 22'b0000000000000000001110, 22'b1111111111111110011001, 22'b1111111111111110101110, 22'b1111111111111111111101, 22'b1111111111111101000101, 22'b1111111111111110110110, 22'b1111111111111101111010, 22'b0000000000000001100000, 22'b0000000000000000110111, 22'b1111111111111010010100, 22'b0000000000000000000001, 22'b1111111111111111111100, 22'b1111111111111111101111, 22'b0000000000000010010000, 22'b1111111111111111010110, 22'b1111111111111111000111, 22'b1111111111111111000100, 22'b1111111111111111111110, 22'b0000000000001000101011, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b1111111111111111101100, 22'b0000000000001010001001, 22'b0000000000000110000010, 22'b0000000000000001000101, 22'b1111111111111100111010, 22'b1111111111111111101011, 22'b0000000000000010000101, 22'b0000000000000001110101}, 
{22'b0000000000000001000101, 22'b0000000000000001010000, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b1111111111110001000000, 22'b0000000000000001011001, 22'b0000000000000000110010, 22'b1111111111111111111111, 22'b0000000000000000000001, 22'b1111111111111010100100, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b1111111111111010110110, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b1111111111110100100111, 22'b0000000000000000010011, 22'b1111111111111111111110, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b0000000000000100001000, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b0000000000001110100101, 22'b0000000000001010111000, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b1111111111111000100001, 22'b0000000000000000000000, 22'b1111111111111111111111}, 
{22'b0000000000000010011011, 22'b0000000000000001101100, 22'b0000000000001000000110, 22'b1111111111111000000011, 22'b0000000000000100001111, 22'b0000000000000011110011, 22'b0000000000000000001100, 22'b0000000000000110001000, 22'b0000000000000000011000, 22'b1111111111111111100111, 22'b0000000000000001001100, 22'b0000000000000000001011, 22'b1111111111111111111110, 22'b0000000000000011110111, 22'b1111111111111111110100, 22'b1111111111111110101110, 22'b0000000000000000000001, 22'b0000000000000001000001, 22'b1111111111111110011101, 22'b0000000000000011001010, 22'b0000000000000001000010, 22'b1111111111101101011011, 22'b1111111111111100010101, 22'b0000000000000010111011, 22'b1111111111111111111111, 22'b1111111111101111110101, 22'b1111111111111011111101, 22'b1111111111111111010000, 22'b1111111111111111111110, 22'b1111111111111110001011, 22'b0000000000000000000000, 22'b1111111111111110101110}, 
{22'b0000000000000000000011, 22'b1111111111111111111111, 22'b1111111111111101000100, 22'b1111111111111010100111, 22'b0000000000000001010101, 22'b0000000000000000000000, 22'b0000000000000011000011, 22'b1111111111111111110100, 22'b0000000000000111111111, 22'b1111111111111111110111, 22'b0000000000000000000000, 22'b1111111111110101000000, 22'b1111111111111111111111, 22'b0000000000000100000001, 22'b1111111111111111111111, 22'b1111111111110111101010, 22'b0000000000000000000000, 22'b1111111111111111101000, 22'b0000000000001000011010, 22'b1111111111111111111111, 22'b1111111111110010000001, 22'b1111111111111111111111, 22'b0000000000001000010000, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b0000000000000100011100, 22'b1111111111111100111111, 22'b0000000000000010001101, 22'b0000000000000000000000, 22'b1111111111111001100011, 22'b0000000000000000000000, 22'b0000000000000000000101}, 
{22'b1111111111111001000101, 22'b0000000000000000000010, 22'b0000000000000000000001, 22'b1111111111111111110011, 22'b0000000000001111110111, 22'b1111111111111100000001, 22'b1111111111111111110100, 22'b1111111111111111110001, 22'b1111111111111110100100, 22'b1111111111111110011000, 22'b0000000000000010000101, 22'b0000000000000100010000, 22'b1111111111111110110100, 22'b0000000000000111111111, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b1111111111110110111010, 22'b1111111111111111111110, 22'b0000000000000000000000, 22'b1111111111111101011100, 22'b0000000000000000000100, 22'b0000000000000001001100, 22'b0000000000000000011011, 22'b1111111111111111101101, 22'b1111111111111110010111, 22'b1111111111111001100000, 22'b1111111111110110100010, 22'b0000000000000000000000, 22'b1111111111111100011000, 22'b0000000000000001010001, 22'b1111111111111111111111, 22'b0000000000000010011010}, 
{22'b1111111111110010110001, 22'b1111111111111010111111, 22'b1111111111111011000000, 22'b0000000000000000000000, 22'b0000000000010010010001, 22'b1111111111111000111000, 22'b0000000000000000000000, 22'b1111111111111110010001, 22'b1111111111110010111000, 22'b0000000000000100011011, 22'b1111111111111111111111, 22'b0000000000010010001001, 22'b0000000000000000000000, 22'b1111111111111110011110, 22'b1111111111111111111111, 22'b0000000000000001000000, 22'b1111111111111111011001, 22'b0000000000000000000000, 22'b1111111111111110100000, 22'b0000000000001111110110, 22'b0000000000000001001111, 22'b1111111111111110101010, 22'b0000000000000011100000, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b1111111111111100111000, 22'b1111111111111110100000, 22'b1111111111110001000001, 22'b1111111111111011011000, 22'b1111111111111111111111, 22'b1111111111111111111101, 22'b1111111111111110000111}, 
{22'b0000000000000111001110, 22'b1111111111100110011010, 22'b1111111111101000110100, 22'b1111111111111010100011, 22'b0000000000010101011010, 22'b1111111111111111111111, 22'b1111111111110100111010, 22'b0000000000001000011110, 22'b0000000000000001111001, 22'b0000000000000000000001, 22'b0000000000000110101010, 22'b1111111111110111010100, 22'b0000000000000000000001, 22'b0000000000000000001000, 22'b1111111111111110111111, 22'b0000000000000000100100, 22'b1111111111111100101011, 22'b1111111111100010100000, 22'b0000000000000101010111, 22'b0000000000001011000010, 22'b0000000000001000011110, 22'b0000000000000000000101, 22'b0000000000000000111011, 22'b1111111111110011000110, 22'b1111111111101011110000, 22'b1111111111111111110101, 22'b1111111111110110011010, 22'b1111111111110001010110, 22'b1111111111111001110000, 22'b1111111111100011111011, 22'b0000000000001101011010, 22'b0000000000001101101111}, 
{22'b0000000000000000000000, 22'b0000000000000000000001, 22'b0000000000000000000100, 22'b0000000000000000000000, 22'b0000000000001000010010, 22'b1111111111111010000001, 22'b0000000000000000100100, 22'b0000000000000010010101, 22'b1111111111110100110101, 22'b0000000000000001001011, 22'b1111111111111111110110, 22'b1111111111111111111110, 22'b1111111111111111111111, 22'b0000000000000111101010, 22'b0000000000000001101010, 22'b0000000000000000101100, 22'b0000000000000001111110, 22'b0000000000001010101010, 22'b1111111111111001000000, 22'b0000000000000000000000, 22'b1111111111111010101111, 22'b1111111111111111111111, 22'b0000000000001010000100, 22'b0000000000000000010000, 22'b1111111111111111111010, 22'b1111111111101110000010, 22'b1111111111111111101101, 22'b1111111111111011000011, 22'b1111111111111110000011, 22'b0000000000000000000111, 22'b0000000000000100010100, 22'b0000000000000011010100}, 
{22'b1111111111111110100111, 22'b0000000000000100010010, 22'b1111111111110110010001, 22'b0000000000000000101010, 22'b0000000000000110001100, 22'b1111111111111110101111, 22'b1111111111111111110110, 22'b0000000000000101001110, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b1111111111111101111010, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b1111111111111110111001, 22'b1111111111111100000110, 22'b1111111111111101111000, 22'b1111111111111110001100, 22'b1111111111111101111111, 22'b1111111111111100011111, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b1111111111111110100100, 22'b1111111111111101110111, 22'b0000000000001100101110, 22'b0000000000000000000000, 22'b1111111111110100011110, 22'b1111111111111111101110, 22'b0000000000000011111100, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b0000000000001000000001, 22'b1111111111111111111111}, 
{22'b1111111111111111111111, 22'b0000000000000000001000, 22'b1111111111111111111111, 22'b1111111111111011000000, 22'b1111111111100100011110, 22'b0000000000000000000001, 22'b0000000000000000000000, 22'b1111111111111111110010, 22'b1111111111101100110100, 22'b0000000000000010100111, 22'b1111111111111100110111, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b1111111111110100001010, 22'b1111111111111110100010, 22'b1111111111111111111111, 22'b0000000000000000000010, 22'b0000000000000000010000, 22'b0000000000000001001010, 22'b0000000000001011000011, 22'b1111111111111100001011, 22'b1111111111110110011011, 22'b0000000000000000000000, 22'b1111111111110111101111, 22'b1111111111111100110101, 22'b1111111111111000100110, 22'b1111111111111111110000, 22'b1111111111111111100110, 22'b1111111111111111011010, 22'b1111111111110000111011, 22'b1111111111111110111010, 22'b0000000000000111110000}, 
{22'b0000000000000011100111, 22'b0000000000000111000000, 22'b1111111111111111111011, 22'b0000000000000101000110, 22'b1111111111111001010000, 22'b1111111111111100000001, 22'b0000000000000011000011, 22'b0000000000000010001100, 22'b1111111111111110011111, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b1111111111110101101111, 22'b1111111111111111111111, 22'b0000000000000100100111, 22'b1111111111111100010101, 22'b0000000000000001000111, 22'b1111111111111111111101, 22'b1111111111111111111101, 22'b0000000000000110101000, 22'b1111111111110101100010, 22'b0000000000001000111111, 22'b0000000000000001100001, 22'b0000000000000000000000, 22'b0000000000000110110001, 22'b0000000000000000000110, 22'b1111111111111110110110, 22'b1111111111110011110100, 22'b1111111111111100011111, 22'b1111111111111010100011, 22'b0000000000000101101011}, 
{22'b0000000000000000000000, 22'b0000000000000000001110, 22'b1111111111110100010010, 22'b1111111111111111111011, 22'b0000000000000110100111, 22'b1111111111111011011110, 22'b1111111111111111100111, 22'b1111111111111111111111, 22'b0000000000000000101001, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b1111111111111001011110, 22'b0000000000000011000100, 22'b0000000000000000001100, 22'b0000000000000000000000, 22'b0000000000000001001100, 22'b1111111111111111111111, 22'b1111111111111011001111, 22'b0000000000000000100100, 22'b0000000000000000000000, 22'b1111111111111110111001, 22'b1111111111111111010011, 22'b0000000000001001011110, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b1111111111110110101000, 22'b1111111111110101100010, 22'b0000000000000111101110, 22'b1111111111111111111101, 22'b1111111111111111111111, 22'b0000000000000000111000, 22'b0000000000001001000010}, 
{22'b1111111111110101000110, 22'b1111111111111111111111, 22'b1111111111111001001100, 22'b0000000000000000001000, 22'b1111111111110100101100, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b1111111111111101111010, 22'b1111111111101110111101, 22'b1111111111111111001011, 22'b0000000000000000000000, 22'b1111111111111111101111, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b1111111111111111101110, 22'b1111111111111110011010, 22'b1111111111111011010001, 22'b1111111111111100111100, 22'b0000000000000010000111, 22'b1111111111111111111011, 22'b1111111111111111001100, 22'b0000000000000000000000, 22'b0000000000001010110001, 22'b1111111111111111111111, 22'b0000000000000100110010, 22'b0000000000000010111011, 22'b1111111111111011100110, 22'b0000000000000110110100, 22'b1111111111111110100010, 22'b0000000000000000000000, 22'b1111111111111111111101, 22'b0000000000010010101000}, 
{22'b1111111111110101111100, 22'b0000000000000000111100, 22'b0000000000000001100111, 22'b1111111111111111000110, 22'b0000000000000111110100, 22'b1111111111110110010101, 22'b1111111111111111110001, 22'b0000000000001000011111, 22'b0000000000000101000110, 22'b0000000000000000010010, 22'b1111111111111111111111, 22'b1111111111111101110011, 22'b1111111111111101001000, 22'b1111111111111101111011, 22'b1111111111111110011010, 22'b0000000000000010111000, 22'b1111111111111111111111, 22'b0000000000000000010000, 22'b0000000000000100100001, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b0000000000000000011110, 22'b0000000000001000000100, 22'b0000000000000001011101, 22'b0000000000000000001101, 22'b1111111111111100100011, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b1111111111111111100011, 22'b1111111111111111100111, 22'b1111111111111111111111, 22'b0000000000000010001010}, 
{22'b1111111111111111111111, 22'b0000000000000000000111, 22'b1111111111111001001101, 22'b1111111111111101100111, 22'b0000000000001001000001, 22'b1111111111111111111111, 22'b1111111111111101100001, 22'b0000000000000111110100, 22'b1111111111111110010011, 22'b0000000000001001010101, 22'b0000000000000010101111, 22'b1111111111111100001001, 22'b0000000000000000000001, 22'b0000000000000000000111, 22'b1111111111111111100001, 22'b0000000000000000101011, 22'b1111111111111101100010, 22'b1111111111110111100100, 22'b0000000000001000111001, 22'b0000000000000100111110, 22'b0000000000010100010011, 22'b0000000000000110011011, 22'b0000000000000111111100, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b0000000000000001110101, 22'b0000000000000010100010, 22'b1111111111110010100011, 22'b1111111111111111111111, 22'b1111111111111111110101, 22'b1111111111111111110010}, 
{22'b0000000000000000000001, 22'b1111111111111101001100, 22'b1111111111111100101011, 22'b0000000000000000000000, 22'b1111111111111000001101, 22'b0000000000000000000000, 22'b0000000000000110001000, 22'b0000000000000011011111, 22'b0000000000000001101100, 22'b1111111111111100110101, 22'b0000000000000000000000, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b1111111111111110101000, 22'b0000000000000110011101, 22'b1111111111111111111111, 22'b1111111111111111111110, 22'b1111111111110110010100, 22'b0000000000000000000000, 22'b1111111111111001110101, 22'b1111111111111111111101, 22'b0000000000000000000000, 22'b1111111111111111110111, 22'b0000000000000000011110, 22'b0000000000000000100011, 22'b0000000000000000111001, 22'b0000000000000100011011, 22'b1111111111111101111010, 22'b1111111111111111110000, 22'b1111111111110001101001, 22'b0000000000000010100001}, 
{22'b0000000000001110001000, 22'b1111111111111111101110, 22'b0000000000000010000111, 22'b1111111111111100101001, 22'b1111111111111101010001, 22'b0000000000000001000100, 22'b0000000000000101001000, 22'b0000000000000000000000, 22'b0000000000010000110111, 22'b0000000000000000000000, 22'b1111111111111111010100, 22'b0000000000000000100110, 22'b0000000000000011000000, 22'b1111111111111111111010, 22'b0000000000000001101101, 22'b0000000000000011010011, 22'b1111111111111111110111, 22'b1111111111110001110000, 22'b1111111111111110001100, 22'b1111111111111111111100, 22'b0000000000000011101110, 22'b0000000000000000000011, 22'b1111111111111111111111, 22'b0000000000000011100110, 22'b0000000000000000100100, 22'b1111111111110111100100, 22'b1111111111111100101101, 22'b0000000000000100001110, 22'b1111111111111111000110, 22'b0000000000001000010000, 22'b1111111111111111111101, 22'b1111111111111010010001}, 
{22'b0000000000000000011010, 22'b0000000000000011010000, 22'b1111111111111111111111, 22'b1111111111111110110000, 22'b1111111111110100101101, 22'b1111111111111111111111, 22'b0000000000000001011110, 22'b1111111111111110100001, 22'b0000000000000101010001, 22'b1111111111111110111010, 22'b1111111111111111111110, 22'b1111111111111110111011, 22'b1111111111111111111111, 22'b1111111111111110110100, 22'b0000000000000000000000, 22'b0000000000001010000001, 22'b0000000000000000000000, 22'b1111111111111111111100, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b0000000000000001000101, 22'b0000000000000100000001, 22'b0000000000000000000000, 22'b0000000000000000001000, 22'b0000000000000001000010, 22'b1111111111111111111110, 22'b0000000000000000000000, 22'b0000000000000000101001, 22'b0000000000000000000011, 22'b0000000000000011000110}, 
{22'b1111111111110110000111, 22'b0000000000000100001010, 22'b0000000000000000100100, 22'b1111111111111100101000, 22'b1111111111110011001110, 22'b1111111111111111011010, 22'b0000000000000010001001, 22'b1111111111110011010010, 22'b0000000000010000010111, 22'b0000000000000010010010, 22'b0000000000000000100000, 22'b0000000000000011000001, 22'b0000000000000001011010, 22'b0000000000000000000001, 22'b0000000000001101000011, 22'b1111111111111101010011, 22'b0000000000000000001010, 22'b0000000000000000000000, 22'b1111111111111111110010, 22'b0000000000000000000111, 22'b1111111111110010001011, 22'b0000000000000000100010, 22'b0000000000000100111001, 22'b0000000000000001001100, 22'b0000000000000001001001, 22'b1111111111101010111111, 22'b1111111111110101000101, 22'b1111111111111000010011, 22'b0000000000000000000101, 22'b1111111111111111111100, 22'b0000000000001010011011, 22'b1111111111111001011100}, 
{22'b1111111111111111100101, 22'b1111111111111001110001, 22'b1111111111111100101100, 22'b1111111111110010111011, 22'b1111111111110111101011, 22'b0000000000001010110000, 22'b0000000000001001111010, 22'b1111111111111010100011, 22'b0000000000000001010101, 22'b1111111111111110110000, 22'b1111111111111100111111, 22'b1111111111110111111101, 22'b0000000000000011010011, 22'b1111111111110110111010, 22'b0000000000000110000010, 22'b1111111111111111111111, 22'b0000000000001010101111, 22'b1111111111111111111111, 22'b1111111111111111110000, 22'b1111111111111011101010, 22'b1111111111111110101010, 22'b1111111111111101111011, 22'b1111111111110111011111, 22'b0000000000000010101000, 22'b1111111111111111111111, 22'b1111111111111111110011, 22'b1111111111111000101100, 22'b0000000000001010000100, 22'b0000000000001000111011, 22'b1111111111111101000110, 22'b1111111111101011110100, 22'b0000000000000100100100}, 
{22'b0000000000000000000000, 22'b1111111111111111001011, 22'b1111111111111111111111, 22'b1111111111111100111000, 22'b0000000000000000111010, 22'b0000000000000000010010, 22'b0000000000000010001110, 22'b0000000000000000001011, 22'b0000000000000011110001, 22'b1111111111111111111110, 22'b0000000000000000000000, 22'b0000000000000011000011, 22'b0000000000000000000011, 22'b0000000000000000011001, 22'b1111111111111011110000, 22'b1111111111111100100011, 22'b0000000000000000000000, 22'b0000000000000101110100, 22'b0000000000000001110100, 22'b0000000000000100000001, 22'b1111111111111111011110, 22'b1111111111111010111000, 22'b1111111111111111111111, 22'b0000000000000010011000, 22'b1111111111111111111111, 22'b0000000000000001000010, 22'b1111111111111111110110, 22'b0000000000000010001010, 22'b0000000000000000000000, 22'b0000000000000010101010, 22'b1111111111110011110110, 22'b1111111111111111111111}, 
{22'b0000000000001001111011, 22'b1111111111111111101101, 22'b0000000000000100110011, 22'b1111111111110110001110, 22'b1111111111111001110100, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b0000000000000000111000, 22'b0000000000000000000100, 22'b1111111111111011111110, 22'b0000000000000000000000, 22'b0000000000000000000100, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b1111111111111011110111, 22'b0000000000000100100100, 22'b1111111111111111111100, 22'b1111111111111111000000, 22'b0000000000000000000000, 22'b0000000000000011110101, 22'b1111111111111001100100, 22'b0000000000000011101101, 22'b0000000000000100011110, 22'b0000000000000100001000, 22'b1111111111111111111111, 22'b0000000000010001101001, 22'b1111111111111011000110, 22'b0000000000001011101000, 22'b1111111111111110010110, 22'b1111111111110100011101, 22'b1111111111111010011100, 22'b0000000000000100011101}, 
{22'b1111111111101110100111, 22'b1111111111111111001001, 22'b1111111111111011000100, 22'b1111111111111111111111, 22'b0000000000001000010110, 22'b1111111111111010010010, 22'b1111111111111110000101, 22'b0000000000000111100111, 22'b0000000000000011000001, 22'b1111111111111000011000, 22'b0000000000000000000000, 22'b1111111111111111000110, 22'b1111111111111111101011, 22'b0000000000000100011001, 22'b1111111111111000001000, 22'b1111111111111111101001, 22'b0000000000000000000000, 22'b1111111111111111111110, 22'b1111111111111111011111, 22'b0000000000000000000000, 22'b1111111111111001111010, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b1111111111110101011111, 22'b0000000000000010001111, 22'b0000000000010011110101, 22'b0000000000001011000100, 22'b1111111111111110110110, 22'b1111111111111010110111, 22'b1111111111110001101001, 22'b0000000000000000000000, 22'b1111111111111110011100}, 
{22'b0000000000000000101011, 22'b0000000000000110110101, 22'b0000000000000000101011, 22'b1111111111111011001010, 22'b0000000000000000001001, 22'b1111111111111111001011, 22'b0000000000000000000000, 22'b0000000000000110101010, 22'b0000000000000110111000, 22'b1111111111111011101110, 22'b0000000000000100011111, 22'b0000000000000000110001, 22'b1111111111111111111111, 22'b1111111111111111100010, 22'b1111111111111010111010, 22'b0000000000001000000110, 22'b1111111111111110101001, 22'b1111111111110101101010, 22'b0000000000000011101010, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b0000000000000011101111, 22'b1111111111111101100111, 22'b1111111111111111110110, 22'b1111111111111110010110, 22'b0000000000000010110100, 22'b1111111111111011100000, 22'b0000000000000100010010, 22'b1111111111110100010111, 22'b0000000000000010100100, 22'b1111111111111111111111, 22'b0000000000000101000000}, 
{22'b1111111111111110101000, 22'b0000000000000000000001, 22'b0000000000000010110110, 22'b0000000000000000000000, 22'b1111111111111110000011, 22'b1111111111111111111010, 22'b0000000000000011010010, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b0000000000000000001010, 22'b0000000000000000000000, 22'b0000000000000000101000, 22'b1111111111111100100110, 22'b0000000000000000010101, 22'b0000000000000011100010, 22'b0000000000000001011111, 22'b0000000000000011011000, 22'b1111111111111111111110, 22'b1111111111111111111101, 22'b0000000000000100000110, 22'b0000000000000111111010, 22'b1111111111111100110111, 22'b0000000000000000000000, 22'b1111111111111111111011, 22'b0000000000000000010111, 22'b1111111111110001001111, 22'b1111111111111111111110, 22'b1111111111111101101111, 22'b1111111111111111111111, 22'b0000000000010010000100, 22'b0000000000000000000000, 22'b1111111111111001011010}, 
{22'b1111111111111111001001, 22'b1111111111111100001011, 22'b1111111111111111101101, 22'b0000000000000000001110, 22'b0000000000000010111001, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b1111111111111111010000, 22'b0000000000000010010000, 22'b1111111111111111101111, 22'b0000000000000000000000, 22'b0000000000000001000000, 22'b0000000000001001011100, 22'b1111111111111100101111, 22'b0000000000000000011001, 22'b1111111111100100110110, 22'b1111111111111111101001, 22'b1111111111111110000100, 22'b0000000000000000010000, 22'b1111111111111110011001, 22'b0000000000000010111100, 22'b1111111111111000110101, 22'b0000000000000011101001, 22'b0000000000000011010111, 22'b1111111111111111100101, 22'b1111111111101001001111, 22'b1111111111111000101011, 22'b1111111111111111010011, 22'b1111111111111111011010, 22'b0000000000001100011111, 22'b1111111111111111110100, 22'b0000000000000100111011}, 
{22'b0000000000000001100000, 22'b0000000000000000000000, 22'b0000000000000101100100, 22'b1111111111111100010111, 22'b1111111111111101110011, 22'b0000000000000111100111, 22'b1111111111111010111000, 22'b0000000000000001110101, 22'b1111111111110110000110, 22'b0000000000000000010001, 22'b0000000000000000100010, 22'b1111111111111101010100, 22'b0000000000000000000001, 22'b0000000000000000000000, 22'b1111111111111001111111, 22'b0000000000001101110101, 22'b1111111111111000000110, 22'b1111111111111111100111, 22'b0000000000000011110011, 22'b1111111111111111111111, 22'b0000000000000010001101, 22'b1111111111110000101010, 22'b0000000000001010000001, 22'b1111111111111111111111, 22'b1111111111111100000010, 22'b0000000000001111100000, 22'b0000000000000100101011, 22'b1111111111111010111100, 22'b1111111111111011101100, 22'b1111111111101110110011, 22'b1111111111111111101011, 22'b0000000000000000100000}, 
{22'b1111111111111111111111, 22'b0000000000000000001101, 22'b1111111111111110111000, 22'b1111111111110111011011, 22'b1111111111111111111111, 22'b1111111111110011011100, 22'b0000000000000000000000, 22'b0000000000001001101101, 22'b0000000000000111110100, 22'b0000000000000000100110, 22'b0000000000000000000000, 22'b1111111111111100011110, 22'b0000000000001010101000, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b0000000000001101111000, 22'b0000000000000000000011, 22'b1111111111111110101110, 22'b1111111111111110010111, 22'b1111111111110101101100, 22'b0000000000000100001101, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b0000000000000001000000, 22'b1111111111111101101110, 22'b1111111111110001010000, 22'b0000000000001000110101, 22'b1111111111110001110011, 22'b0000000000000001101000, 22'b1111111111111101011110, 22'b0000000000000000000000}, 
{22'b0000000000000001111101, 22'b0000000000000101111101, 22'b0000000000000000010011, 22'b1111111111111111111001, 22'b1111111111110001010011, 22'b0000000000000000000001, 22'b1111111111111111111111, 22'b0000000000000111110000, 22'b0000000000001000110111, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b1111111111111111111101, 22'b0000000000000000000000, 22'b0000000000000000000100, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b1111111111111111111110, 22'b0000000000000101011100, 22'b1111111111111100101101, 22'b1111111111110010001011, 22'b1111111111111110111100, 22'b1111111111111100110101, 22'b1111111111111100111111, 22'b1111111111111101110010, 22'b1111111111111111111110, 22'b1111111111111101111111, 22'b1111111111111111010011, 22'b1111111111111111101010, 22'b0000000000000100100001, 22'b1111111111111111111111, 22'b0000000000001110110101}
};

localparam logic signed [21:0] bias [32] = '{
22'b0000000000101111001011,  // 1.474280834197998
22'b0000000000010110001000,  // 0.6914801001548767
22'b0000000000101110000110,  // 1.4406442642211914
22'b0000000000101101000011,  // 1.408045768737793
22'b0000000000011111100100,  // 0.9864811301231384
22'b0000000000011011101000,  // 0.8636202812194824
22'b1111111111101100010011,  // -0.6153604388237
22'b0000000000001111011111,  // 0.4839226007461548
22'b0000000000001111100011,  // 0.4862793982028961
22'b0000000000001011111001,  // 0.37162142992019653
22'b0000000000001110101101,  // 0.45989668369293213
22'b0000000000101001100110,  // 1.2998151779174805
22'b1111111111011111011110,  // -1.016528844833374
22'b1111111111110100101110,  // -0.35249894857406616
22'b0000000000001110010001,  // 0.44582197070121765
22'b1111111111111100011010,  // -0.1119980737566948
22'b1111111111111101110110,  // -0.06717441976070404
22'b0000000000000000001001,  // 0.00487547367811203
22'b0000000000000110001110,  // 0.1946917623281479
22'b1111111111100111000011,  // -0.7796769738197327
22'b0000000000010111010100,  // 0.7287401556968689
22'b0000000000110110111000,  // 1.714877724647522
22'b1111111111001100111001,  // -1.5971007347106934
22'b0000000000000010010111,  // 0.07393483817577362
22'b0000000000001010010100,  // 0.3225609362125397
22'b0000000000011011000011,  // 0.8453295230865479
22'b0000000000011100110000,  // 0.898597240447998
22'b0000000000001000001001,  // 0.2548799514770508
22'b0000000000011111001001,  // 0.9735668301582336
22'b0000000000100100000010,  // 1.1261906623840332
22'b0000000000001110010100,  // 0.44768181443214417
22'b1111111110110100001111   // -2.3676068782806396
};
endpackage