//Width: 37
//Int: 13
package dense_4_gen;

localparam logic signed [36:0] weights [32][5] = '{
{37'b1111111111111111111001111010110111010, 37'b0000000000000010100001100110011001000, 37'b1111111111111101100111011100001100111, 37'b0000000000000000100001101100111000111, 37'b1111111111111111001001100101111111000},
{37'b1111111111111011100010011110010100011, 37'b1111111111111111100011110111100100001, 37'b0000000000000011101011101001111110100, 37'b1111111111111111111001101101000110101, 37'b0000000000000000001000100100000011111},
{37'b0000000000000010111110001111010111010, 37'b0000000000000001101100011010001100001, 37'b1111111111111111110001101011101110111, 37'b1111111111111100110000011101000001111, 37'b1111111111111110010100000011101111111},
{37'b1111111111111100111111101101000110001, 37'b1111111111111101000001000100101110001, 37'b1111111111111111000110110001101101100, 37'b0000000000000010011101100111100000010, 37'b0000000000000001111000010101000010000},
{37'b0000000000000000111110100011111011011, 37'b0000000000000001000001111000011110010, 37'b0000000000000001010000011011101111011, 37'b1111111111111111110110101000001011111, 37'b1111111111110111111001011000111011000},
{37'b0000000000000010100111011100101010010, 37'b1111111111111100110110000100001000110, 37'b0000000000000001011100111001000111110, 37'b1111111111111110101101011101011001101, 37'b1111111111111110101000110011010011101},
{37'b1111111111111100110010100010000110000, 37'b0000000000000000010010001110010101011, 37'b1111111111111111111111111111100111011, 37'b0000000000000001011001001010101011100, 37'b0000000000000000100011010101111100100},
{37'b1111111111111111111111000001001111101, 37'b0000000000000010010001101010011001000, 37'b1111111111111100110111010111111111011, 37'b0000000000000001010011010011100101000, 37'b0000000000000001000101101100011110110},
{37'b0000000000000001010011101000000101100, 37'b1111111111111110101001010001110010100, 37'b0000000000000000000000101010010101110, 37'b1111111111111100010011101110111010101, 37'b1111111111111110000000101011001011010},
{37'b1111111111111111111111111000101010011, 37'b1111111111111101110111101010110010111, 37'b0000000000000001011011000100011100010, 37'b0000000000000011011100001000010001101, 37'b0000000000000000000000000000101101001},
{37'b1111111111111110111101011100001101101, 37'b1111111111111110110101111111011001001, 37'b0000000000000000000000000000010100000, 37'b0000000000000100101001101011011000111, 37'b1111111111111101110110111101111000001},
{37'b0000000000000001010110101110111100010, 37'b0000000000000001110101010101101100110, 37'b1111111111111101010001111000011110111, 37'b1111111111111111110001111010000101000, 37'b0000000000000000111110010101010010101},
{37'b0000000000000000000000000010011100110, 37'b0000000000000001010101110101001101100, 37'b0000000000000000000100100101001011111, 37'b1111111111111110010101100110011100001, 37'b1111111111111011000001000110011000111},
{37'b0000000000000001011010110000011001000, 37'b0000000000000000100000101011000110010, 37'b0000000000000011010110110011111011110, 37'b1111111111111111011100001001001001111, 37'b1111111111111100100100111101111001101},
{37'b0000000000000000101110011111001101100, 37'b1111111111111111100111010110011111001, 37'b1111111111111101000111011100101110010, 37'b1111111111111111101111000110110011111, 37'b0000000000000100010010100110101001100},
{37'b1111111111111100001101010000100111101, 37'b1111111111111110000010111010111110111, 37'b1111111111111110001110000111011101001, 37'b0000000000000011001100001110011001000, 37'b0000000000000000010000011011100011100},
{37'b0000000000000010110001000011010000011, 37'b1111111111111110101000000100001010101, 37'b1111111111111110111010100001010000101, 37'b1111111111111110001100011111110011111, 37'b1111111111111111100001010101000100110},
{37'b0000000000000001100011110110100000100, 37'b1111111111111111101011010001010101111, 37'b1111111111111100101100111001111001011, 37'b1111111111111111110000010100010001011, 37'b0000000000000000100100001100000100110},
{37'b0000000000000010000100010110010111000, 37'b0000000000000000010101010010100110000, 37'b1111111111111110010000011000011010011, 37'b0000000000000000000000000000010100110, 37'b1111111111111100111111100111111011000},
{37'b0000000000000001110110011111010110000, 37'b1111111111111111010011101100011111001, 37'b1111111111111110010011000011101010010, 37'b0000000000000001101010000101110010011, 37'b0000000000000000110000101100001100001},
{37'b0000000000000000100010101011100010111, 37'b1111111111111111110000011111010001010, 37'b0000000000000010011000010111111011110, 37'b1111111111111100100011010110011100101, 37'b1111111111111111110101000110101100001},
{37'b0000000000000000000000000000000000011, 37'b0000000000000000111100010111000001001, 37'b0000000000000011111001001000110000010, 37'b1111111111111011110110101001110110110, 37'b1111111111111011000011110010010010010},
{37'b1111111111111111001101101111101111010, 37'b0000000000000000111000001011000000000, 37'b0000000000000001011010101100111000100, 37'b1111111111111101001001010010001100001, 37'b0000000000000100001011011100101001001},
{37'b1111111111111111111111110011101000110, 37'b0000000000000001010100011010111011101, 37'b0000000000000010010000101110110101100, 37'b0000000000000000010011011100011011011, 37'b1111111111111011011011000111011111110},
{37'b1111111111111110101001010100101110111, 37'b0000000000000010111010100001111011101, 37'b1111111111111110001101100001000011110, 37'b0000000000000000000010111011011101111, 37'b0000000000000011000110101111000110000},
{37'b0000000000000000001101011101001111001, 37'b0000000000000010001000000001011110010, 37'b0000000000000000001111001000101001000, 37'b1111111111111010000001000011000111100, 37'b0000000000000100011000101100011000010},
{37'b1111111111111100010100101001110011011, 37'b1111111111111110000011010011010110010, 37'b0000000000000001101101101000011101110, 37'b0000000000000001111101001100101101011, 37'b0000000000000001100111010011100010001},
{37'b0000000000000000000010000100101000010, 37'b0000000000000001111011011010110100110, 37'b1111111111111111101101010011100001100, 37'b1111111111111110110010111100101011010, 37'b0000000000000000010000001100010000010},
{37'b1111111111111111001010101001001001110, 37'b0000000000000001111110000010011000100, 37'b1111111111111011111110000000011111001, 37'b0000000000000001000111000011001011110, 37'b1111111111111110101110111011100010111},
{37'b1111111111111111110110100111001101111, 37'b0000000000000001001000010000000110011, 37'b1111111111111110101001100111011100011, 37'b1111111111111100110010111110001110110, 37'b0000000000000100101111111001111100110},
{37'b0000000000000011100101110101110000001, 37'b0000000000000000100011110011001110000, 37'b0000000000000010100110001001011110110, 37'b1111111111111011010010000001101001001, 37'b1111111111111101011110101001110001111},
{37'b1111111111111111100001101100110100001, 37'b1111111111111100111010010011000011111, 37'b0000000000000010111011010010000110100, 37'b0000000000000000100100010000110010111, 37'b0000000000000001000001010010011001111}
};
localparam logic signed [36:0] bias [5] = '{
37'b1111111111111111100000001000110011010,
37'b1111111111111111011111111001010000111,
37'b1111111111111111011100000101100010110,
37'b0000000000000000101010000001100001000,
37'b0000000000000001101110010111111011111
};
endpackage