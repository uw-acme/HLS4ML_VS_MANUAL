// Width: 13
// NFRAC: 6
package dense_1_13_6;

localparam logic signed [12:0] weights [16][64] = '{ 
{13'b0000000010000, 13'b1111111010110, 13'b1111111110100, 13'b1111111110001, 13'b1111111100110, 13'b0000000000111, 13'b1111110111101, 13'b0000000000000, 13'b0000000000011, 13'b0000000010000, 13'b0000000000000, 13'b1111111100110, 13'b1111111111111, 13'b0000000001101, 13'b0000000000010, 13'b1111111101111, 13'b0000000001110, 13'b0000000000011, 13'b0000000000000, 13'b1111111111111, 13'b0000000011000, 13'b1111111101010, 13'b1111111111110, 13'b0000000011110, 13'b1111111101011, 13'b1111111010100, 13'b1111111101110, 13'b1111111110011, 13'b1111111111001, 13'b1111111111111, 13'b0000000000010, 13'b0000000001111, 13'b0000000001100, 13'b1111111111111, 13'b0000000000000, 13'b0000000010011, 13'b1111111111110, 13'b1111111101111, 13'b0000000000001, 13'b0000000001100, 13'b1111111111111, 13'b0000000010001, 13'b1111111101110, 13'b0000000111011, 13'b1111111111111, 13'b0000000011100, 13'b0000000000000, 13'b0000000001011, 13'b0000000001100, 13'b1111111111110, 13'b0000000000000, 13'b0000000001010, 13'b0000000001101, 13'b0000000000100, 13'b1111111111000, 13'b1111111101100, 13'b0000000100010, 13'b1111111100000, 13'b0000000011101, 13'b1111111101001, 13'b0000000110010, 13'b1111111111111, 13'b0000000000000, 13'b0000000000101}, 
{13'b0000000000000, 13'b1111111101011, 13'b1111111110111, 13'b1111111101110, 13'b1111111101011, 13'b0000000000110, 13'b1111111001111, 13'b1111111111111, 13'b1111111110001, 13'b0000000001011, 13'b0000000000000, 13'b1111111111010, 13'b0000000001100, 13'b0000000000000, 13'b1111111111111, 13'b0000000001101, 13'b1111111111111, 13'b0000000000000, 13'b1111111110100, 13'b1111111101111, 13'b0000000011100, 13'b1111111111010, 13'b0000000000011, 13'b0000000101100, 13'b0000000010000, 13'b1111111110001, 13'b1111111110001, 13'b1111111111111, 13'b1111111111001, 13'b1111111100110, 13'b1111111111100, 13'b0000000011101, 13'b0000000010001, 13'b0000000100011, 13'b0000000101000, 13'b0000000000011, 13'b1111111111000, 13'b1111111100100, 13'b0000000000011, 13'b0000000001100, 13'b0000000000001, 13'b0000000001101, 13'b1111111110010, 13'b0000000010000, 13'b0000000001011, 13'b0000000000011, 13'b1111111101010, 13'b0000000000101, 13'b0000000010000, 13'b0000000000001, 13'b0000000000001, 13'b0000001001010, 13'b1111111111011, 13'b1111111111001, 13'b1111111111100, 13'b1111111111111, 13'b0000000010000, 13'b1111111101000, 13'b0000000111111, 13'b0000000000000, 13'b0000000100001, 13'b0000000001111, 13'b0000000110100, 13'b0000000001001}, 
{13'b1111111111111, 13'b0000000000000, 13'b1111111111010, 13'b1111111110100, 13'b1111111110100, 13'b0000000000010, 13'b0000001011110, 13'b1111111111111, 13'b1111110101110, 13'b1111111111111, 13'b1111111111111, 13'b1111111111110, 13'b1111111110001, 13'b0000000000000, 13'b1111111111111, 13'b0000000001010, 13'b0000000111001, 13'b1111111111111, 13'b0000000000100, 13'b0000000000000, 13'b0000000011010, 13'b1111111010001, 13'b0000000100100, 13'b1111111010010, 13'b0000000111100, 13'b1111111101001, 13'b1111111110000, 13'b1111111010010, 13'b0000001010001, 13'b0000000010001, 13'b0000000000000, 13'b0000000100001, 13'b0000001000001, 13'b1111110110011, 13'b1111111111001, 13'b0000000000010, 13'b1111111110001, 13'b0000000111001, 13'b1111111111101, 13'b0000000010100, 13'b0000000010101, 13'b0000000010111, 13'b1111111111111, 13'b1111111111111, 13'b1111111111110, 13'b0000000001010, 13'b1111111101110, 13'b1111111110101, 13'b1111111111110, 13'b0000000011001, 13'b1111111110100, 13'b0000000001001, 13'b1111111111111, 13'b0000000001000, 13'b1111111110100, 13'b1111111111111, 13'b1111111101100, 13'b1111111010101, 13'b1111111111111, 13'b0000000000000, 13'b0000001100010, 13'b0000000000000, 13'b1111111111111, 13'b1111111101100}, 
{13'b1111111100010, 13'b1111111101000, 13'b1111111010011, 13'b0000000010011, 13'b1111111101011, 13'b1111110101001, 13'b1111111111000, 13'b1111111101100, 13'b0000000001110, 13'b1111111111111, 13'b0000001010000, 13'b1111111111001, 13'b1111111001101, 13'b0000000100101, 13'b0000000000001, 13'b1111111111111, 13'b1111111100011, 13'b1111111111111, 13'b0000000000000, 13'b1111111110001, 13'b1111110110110, 13'b1111111111000, 13'b1111111010011, 13'b0000000001100, 13'b1111111100111, 13'b1111111000101, 13'b0000000010100, 13'b0000000101111, 13'b0000001010010, 13'b1111111100010, 13'b1111111011010, 13'b0000000000100, 13'b0000000100000, 13'b1111111001010, 13'b1111111101011, 13'b0000000000000, 13'b1111111010001, 13'b0000000001111, 13'b1111111100011, 13'b0000000000111, 13'b0000000011101, 13'b0000000001010, 13'b0000000000000, 13'b0000000000001, 13'b0000000100011, 13'b1111111110011, 13'b1111111111111, 13'b1111111101001, 13'b1111111111111, 13'b1111111111001, 13'b1111111011000, 13'b0000000000101, 13'b1111111111111, 13'b0000000001101, 13'b0000000010100, 13'b0000000101001, 13'b1111111000010, 13'b1111111000100, 13'b1111111010010, 13'b0000000110111, 13'b0000001101111, 13'b1111111000110, 13'b1111111111100, 13'b0000000011011}, 
{13'b0000000010101, 13'b1111111011000, 13'b1111111101111, 13'b1111111111111, 13'b1111111110110, 13'b0000000010101, 13'b0000000001100, 13'b1111111111111, 13'b1111111011001, 13'b1111111110000, 13'b1111111101000, 13'b0000000000011, 13'b0000000000000, 13'b0000000000000, 13'b1111111111101, 13'b0000000010110, 13'b0000000001000, 13'b1111111100110, 13'b0000000000001, 13'b0000000000000, 13'b0000000001101, 13'b1111111111000, 13'b0000000000100, 13'b1111111111110, 13'b0000001000100, 13'b1111111110100, 13'b1111111101110, 13'b1111111100110, 13'b0000000000000, 13'b0000000001010, 13'b0000000000111, 13'b0000000010001, 13'b1111111111111, 13'b0000000000100, 13'b0000000001000, 13'b1111111111111, 13'b0000000000000, 13'b0000000111000, 13'b1111111101101, 13'b1111111111011, 13'b0000000011011, 13'b0000000001111, 13'b1111111100000, 13'b0000000000000, 13'b1111110111011, 13'b1111111111111, 13'b1111111111000, 13'b0000000000000, 13'b1111111111111, 13'b1111111111110, 13'b1111111111111, 13'b0000000001100, 13'b1111111111111, 13'b0000000010100, 13'b1111111110011, 13'b1111111010000, 13'b1111111100010, 13'b1111111011111, 13'b1111111011000, 13'b0000000101111, 13'b0000001010111, 13'b0000000110010, 13'b0000000000111, 13'b1111111111111}, 
{13'b1111111100011, 13'b1111111010111, 13'b0000000000000, 13'b0000000010011, 13'b0000000010010, 13'b1111111110010, 13'b0000000100101, 13'b1111111111111, 13'b0000000001111, 13'b1111111111111, 13'b1111111111111, 13'b1111111111011, 13'b1111111110100, 13'b0000000100101, 13'b1111111111010, 13'b0000000000000, 13'b1111111011000, 13'b1111111101001, 13'b0000000000000, 13'b1111111111111, 13'b1111111111100, 13'b1111111101011, 13'b1111111101011, 13'b0000000011101, 13'b1111111101011, 13'b1111111111111, 13'b0000000010000, 13'b1111111111011, 13'b1111111000100, 13'b1111111111111, 13'b1111111111011, 13'b1111111111111, 13'b1111111111111, 13'b0000000000010, 13'b0000000001000, 13'b0000000010110, 13'b0000000000000, 13'b1111111111001, 13'b1111111101111, 13'b1111111111111, 13'b1111111110101, 13'b1111111011110, 13'b0000000011001, 13'b0000000000000, 13'b0000000100110, 13'b0000000000000, 13'b1111111111111, 13'b0000000000110, 13'b1111111100101, 13'b0000000001110, 13'b0000000000000, 13'b1111111111001, 13'b1111111101000, 13'b0000000011000, 13'b1111111111111, 13'b0000000010110, 13'b0000000001101, 13'b0000000001101, 13'b1111111111110, 13'b1111111111111, 13'b1111111001100, 13'b1111111110111, 13'b1111111111100, 13'b1111111111111}, 
{13'b1111111101101, 13'b1111111101010, 13'b1111111100100, 13'b1111111111011, 13'b1111111110111, 13'b0000000000110, 13'b1111111010011, 13'b1111111110110, 13'b1111111110001, 13'b1111111111111, 13'b1111111101101, 13'b0000000010110, 13'b0000000000010, 13'b0000000001000, 13'b0000000010011, 13'b0000000000000, 13'b0000000110011, 13'b0000000000101, 13'b0000000001111, 13'b0000000010001, 13'b1111111110101, 13'b0000000010111, 13'b1111111110000, 13'b1111111011111, 13'b0000000001011, 13'b0000000100001, 13'b1111111111111, 13'b0000000000011, 13'b1111111000011, 13'b0000000010010, 13'b0000000010001, 13'b1111111101000, 13'b0000000011110, 13'b0000000101010, 13'b0000000000000, 13'b0000000010101, 13'b1111111111111, 13'b0000000010010, 13'b0000000001100, 13'b0000000000000, 13'b1111111111000, 13'b1111111101000, 13'b0000000001001, 13'b0000000011110, 13'b0000000100001, 13'b1111111110101, 13'b1111111111010, 13'b1111111110011, 13'b1111111110111, 13'b0000000000111, 13'b0000000000000, 13'b0000000000010, 13'b0000000000000, 13'b0000000001011, 13'b1111111110100, 13'b0000000110001, 13'b0000000010110, 13'b1111111111110, 13'b0000000011000, 13'b0000000001101, 13'b1111110010111, 13'b1111111011011, 13'b1111111110100, 13'b1111111111111}, 
{13'b0000000000000, 13'b0000000001111, 13'b1111111111111, 13'b1111111111111, 13'b1111111101011, 13'b1111111111110, 13'b1111111101111, 13'b0000000000000, 13'b0000000000001, 13'b0000000011000, 13'b0000000000000, 13'b1111111100111, 13'b1111111111011, 13'b0000000000000, 13'b1111111111100, 13'b1111111100011, 13'b1111111001001, 13'b1111111111111, 13'b1111111011001, 13'b1111111100011, 13'b1111111100111, 13'b0000000010110, 13'b0000000000011, 13'b1111111110110, 13'b1111111100100, 13'b0000000001001, 13'b0000000000000, 13'b0000000011111, 13'b0000000110011, 13'b1111111111101, 13'b0000000000000, 13'b0000000001110, 13'b1111111010100, 13'b1111111101000, 13'b0000000000011, 13'b0000000000101, 13'b1111111101110, 13'b0000000001111, 13'b0000000001000, 13'b1111111110110, 13'b1111111100101, 13'b1111111111101, 13'b0000000000010, 13'b1111111110101, 13'b0000000000011, 13'b0000000001110, 13'b1111111111000, 13'b0000000000001, 13'b0000000000000, 13'b1111111110010, 13'b1111111100111, 13'b0000000011010, 13'b0000000001000, 13'b1111111110100, 13'b0000000001000, 13'b1111111111100, 13'b1111111100001, 13'b1111111110111, 13'b1111111111100, 13'b1111111111011, 13'b0000000110101, 13'b0000000001100, 13'b1111111111100, 13'b1111111111111}, 
{13'b0000000000000, 13'b0000000100101, 13'b1111111011010, 13'b1111111110001, 13'b0000000010100, 13'b1111111110010, 13'b0000001001101, 13'b1111111101101, 13'b1111111111111, 13'b0000000010010, 13'b0000000010000, 13'b1111111111111, 13'b1111111111100, 13'b1111111100001, 13'b0000000010010, 13'b0000000001010, 13'b1111111110011, 13'b1111111111111, 13'b0000000000000, 13'b0000000000000, 13'b0000000010000, 13'b1111111100010, 13'b0000000011001, 13'b0000000100111, 13'b1111111111010, 13'b1111111111111, 13'b1111111111110, 13'b1111111111111, 13'b0000000101111, 13'b0000000000000, 13'b1111111101110, 13'b0000000000000, 13'b0000000011000, 13'b1111111001100, 13'b1111111011101, 13'b0000000001100, 13'b0000000001000, 13'b1111111011011, 13'b1111111110011, 13'b1111111110010, 13'b0000000011001, 13'b0000000011001, 13'b0000000000000, 13'b1111111101110, 13'b0000000000000, 13'b0000000011001, 13'b1111111111100, 13'b1111111111111, 13'b0000000000000, 13'b0000000001111, 13'b1111111111100, 13'b1111111110011, 13'b0000000010110, 13'b1111111110010, 13'b0000000010001, 13'b0000000100101, 13'b0000000000010, 13'b0000000010000, 13'b1111111100110, 13'b1111111101000, 13'b0000000110101, 13'b1111111110111, 13'b0000000000010, 13'b1111111111010}, 
{13'b0000000000001, 13'b1111111100011, 13'b0000000010111, 13'b1111111101101, 13'b1111111111111, 13'b0000000001101, 13'b1111111011010, 13'b0000000001100, 13'b0000000011111, 13'b0000000001001, 13'b0000000010111, 13'b0000000010100, 13'b1111111101100, 13'b1111111111011, 13'b1111111111100, 13'b0000000000000, 13'b1111111000010, 13'b0000000010100, 13'b1111111111101, 13'b0000000000001, 13'b1111111101001, 13'b0000000000100, 13'b0000000001001, 13'b1111111111111, 13'b1111111100010, 13'b1111111111100, 13'b1111111111010, 13'b0000001001111, 13'b1111111010101, 13'b0000000000100, 13'b0000000000110, 13'b1111111111100, 13'b1111111110001, 13'b0000000000111, 13'b1111111111010, 13'b1111111110111, 13'b1111111110100, 13'b1111111110010, 13'b1111111111110, 13'b1111111101100, 13'b0000000010100, 13'b0000000000111, 13'b0000000011111, 13'b0000000000101, 13'b0000000000010, 13'b1111111101101, 13'b0000000000000, 13'b1111111111111, 13'b1111111111111, 13'b0000000001100, 13'b0000000001011, 13'b0000000010010, 13'b1111111111111, 13'b1111111101101, 13'b0000000000000, 13'b0000000000000, 13'b0000000010100, 13'b1111111110011, 13'b1111111011100, 13'b0000000100011, 13'b1111111101101, 13'b0000001001010, 13'b1111111111110, 13'b1111111101001}, 
{13'b1111111011011, 13'b1111111111111, 13'b1111111100101, 13'b0000000001110, 13'b0000000010000, 13'b1111111111001, 13'b0000000100001, 13'b1111111110101, 13'b1111111100001, 13'b1111111101000, 13'b1111111101111, 13'b1111111100001, 13'b1111111110001, 13'b0000000001100, 13'b0000000000000, 13'b0000000000000, 13'b0000000110101, 13'b1111111111101, 13'b1111111111111, 13'b0000000011010, 13'b0000000010010, 13'b1111111011010, 13'b1111111100111, 13'b0000000001100, 13'b1111111100100, 13'b1111111111110, 13'b1111111101111, 13'b1111111101010, 13'b1111111100100, 13'b0000000010011, 13'b0000000001110, 13'b1111111110110, 13'b1111111111011, 13'b1111111000001, 13'b1111111110100, 13'b0000000000011, 13'b1111111110111, 13'b1111111101101, 13'b1111111111111, 13'b0000000000111, 13'b1111111111000, 13'b1111111111111, 13'b1111111111101, 13'b1111111010101, 13'b0000000000000, 13'b0000000000000, 13'b0000000010101, 13'b1111111111000, 13'b0000000011011, 13'b1111111110011, 13'b0000000010010, 13'b1111111111111, 13'b0000000001110, 13'b1111111100110, 13'b1111111111111, 13'b0000000100000, 13'b0000000010100, 13'b0000000010010, 13'b0000000000001, 13'b1111111100110, 13'b1111111101100, 13'b1111111010100, 13'b1111111111111, 13'b0000000000110}, 
{13'b0000000010011, 13'b0000000000000, 13'b0000000001000, 13'b1111111111111, 13'b0000000001001, 13'b1111111110111, 13'b0000000001111, 13'b0000000000010, 13'b0000000001000, 13'b0000000010101, 13'b1111111101111, 13'b1111111111110, 13'b1111111111111, 13'b1111111111111, 13'b1111111010101, 13'b1111111101100, 13'b0000000101000, 13'b1111111111110, 13'b1111111111100, 13'b0000000000000, 13'b1111111100111, 13'b0000000000000, 13'b0000000010000, 13'b0000000000010, 13'b0000000000010, 13'b0000000010101, 13'b0000000000000, 13'b0000000000010, 13'b0000000000000, 13'b1111111111100, 13'b1111111110011, 13'b1111111010101, 13'b0000000010000, 13'b0000000010101, 13'b1111111111110, 13'b1111111110000, 13'b0000000000000, 13'b1111111010110, 13'b1111111111101, 13'b1111111111111, 13'b0000000001100, 13'b1111111110111, 13'b1111111111111, 13'b0000000110110, 13'b0000000011100, 13'b1111111111111, 13'b1111111111111, 13'b1111111111111, 13'b1111111110000, 13'b0000000001001, 13'b0000000001001, 13'b0000000001011, 13'b0000000001010, 13'b0000000011000, 13'b0000000010110, 13'b0000000101010, 13'b1111111110111, 13'b0000000011001, 13'b0000000001001, 13'b1111111101011, 13'b0000000000111, 13'b1111111100111, 13'b1111111100011, 13'b1111111100000}, 
{13'b0000000000000, 13'b0000000001110, 13'b1111111110011, 13'b0000000000000, 13'b1111111111100, 13'b1111111111101, 13'b1111111010101, 13'b1111111111111, 13'b0000000010000, 13'b0000000001111, 13'b0000000001111, 13'b1111111100110, 13'b1111111111010, 13'b0000000010010, 13'b1111111111111, 13'b0000000000000, 13'b1111111001010, 13'b1111111111111, 13'b0000000010111, 13'b0000000000100, 13'b0000000001111, 13'b1111111111000, 13'b0000000001111, 13'b0000000011001, 13'b1111111101001, 13'b1111111101110, 13'b1111111111111, 13'b1111111111010, 13'b0000000000100, 13'b0000000000000, 13'b1111111111111, 13'b0000000010100, 13'b1111111010000, 13'b0000000010111, 13'b0000000100000, 13'b0000000000111, 13'b0000000000111, 13'b1111111111001, 13'b0000000000111, 13'b1111111111001, 13'b1111111101111, 13'b1111111111100, 13'b0000000001010, 13'b0000000101100, 13'b1111111001001, 13'b1111111100011, 13'b0000000001100, 13'b1111111111001, 13'b0000000011100, 13'b1111111110000, 13'b1111111101010, 13'b1111111101110, 13'b1111111111111, 13'b0000000000111, 13'b1111111110101, 13'b1111111001010, 13'b1111111110110, 13'b1111111111111, 13'b0000000000010, 13'b1111111011000, 13'b0000001000111, 13'b1111111011101, 13'b0000000100010, 13'b0000000001001}, 
{13'b0000000000101, 13'b1111111110011, 13'b0000000101000, 13'b1111111101100, 13'b1111111100010, 13'b0000000000101, 13'b0000000010011, 13'b0000000010011, 13'b1111111110100, 13'b1111111110101, 13'b0000000000011, 13'b0000000001110, 13'b0000000001111, 13'b0000000000011, 13'b1111111110010, 13'b0000000001000, 13'b0000000011110, 13'b1111111111111, 13'b1111111101110, 13'b0000000000000, 13'b0000000000100, 13'b0000000000001, 13'b1111111101101, 13'b0000000000111, 13'b0000000110010, 13'b0000000000000, 13'b0000000001011, 13'b1111111001101, 13'b1111111111011, 13'b0000000000000, 13'b1111111110011, 13'b1111111101100, 13'b0000000011101, 13'b1111111111110, 13'b1111111111101, 13'b1111111101100, 13'b0000000001000, 13'b0000000010010, 13'b1111111111111, 13'b1111111111101, 13'b1111111110100, 13'b0000000001110, 13'b0000000000000, 13'b1111111010100, 13'b0000000010011, 13'b0000000011001, 13'b1111111111111, 13'b0000000000001, 13'b1111111100100, 13'b1111111111011, 13'b1111111111111, 13'b1111111101011, 13'b0000000000000, 13'b1111111110100, 13'b0000000000011, 13'b1111111001011, 13'b1111111111111, 13'b1111111111111, 13'b0000000010001, 13'b0000000100100, 13'b1111111010011, 13'b0000000100001, 13'b0000000000010, 13'b1111111111011}, 
{13'b0000000010010, 13'b0000001001111, 13'b0000000011111, 13'b0000000010010, 13'b1111111100001, 13'b1111111101011, 13'b1111101011001, 13'b1111111100010, 13'b0000000011001, 13'b1111111111111, 13'b0000000010010, 13'b0000000110111, 13'b0000000000100, 13'b0000000000000, 13'b1111111111110, 13'b0000000000000, 13'b1111111110011, 13'b1111111110011, 13'b0000000001110, 13'b1111111011111, 13'b1111111010101, 13'b1111111111001, 13'b1111111011010, 13'b0000000000001, 13'b1111101101110, 13'b0000000110100, 13'b0000000111111, 13'b0000000100110, 13'b1111110010000, 13'b1111111101011, 13'b1111111010011, 13'b1111111001010, 13'b1111101011110, 13'b0000000101011, 13'b1111111111101, 13'b0000000010100, 13'b0000000000001, 13'b1111110100100, 13'b0000000000000, 13'b0000000000000, 13'b0000000000010, 13'b0000001000001, 13'b1111111110010, 13'b1111111010110, 13'b0000000111001, 13'b1111111100011, 13'b1111111101011, 13'b1111111100110, 13'b0000000011110, 13'b0000000100010, 13'b1111111111011, 13'b1111111101001, 13'b1111111111111, 13'b1111111111000, 13'b0000000000000, 13'b1111111100111, 13'b0000000100110, 13'b0000001000101, 13'b0000000101101, 13'b1111111000101, 13'b1111100010011, 13'b0000000111000, 13'b0000000000101, 13'b0000000010100}, 
{13'b1111111110000, 13'b0000000010101, 13'b0000000010100, 13'b1111111111111, 13'b1111111101000, 13'b1111111111010, 13'b1111111100111, 13'b1111111111100, 13'b0000000001001, 13'b1111111111011, 13'b1111111111110, 13'b1111111111101, 13'b1111111111111, 13'b1111111110100, 13'b1111111111110, 13'b1111111111001, 13'b0000000010100, 13'b1111111111111, 13'b1111111010110, 13'b0000000011101, 13'b0000000100110, 13'b0000000011010, 13'b1111111101011, 13'b1111111110111, 13'b1111111101001, 13'b1111111101101, 13'b0000000001110, 13'b0000000001110, 13'b0000000001110, 13'b0000000010111, 13'b0000000000010, 13'b0000000011000, 13'b1111111111101, 13'b0000000000000, 13'b0000000010011, 13'b0000000001000, 13'b1111111111011, 13'b1111111111111, 13'b0000000000000, 13'b1111111101101, 13'b1111111110001, 13'b1111111111000, 13'b1111111101001, 13'b0000000011100, 13'b0000000000000, 13'b1111111111111, 13'b1111111111010, 13'b1111111110110, 13'b1111111001100, 13'b1111111111101, 13'b1111111110001, 13'b1111111110110, 13'b1111111111001, 13'b0000000010000, 13'b0000000101011, 13'b0000000001011, 13'b1111111111111, 13'b1111111101010, 13'b1111111111110, 13'b0000000000000, 13'b0000000010100, 13'b1111111111110, 13'b0000000000010, 13'b0000000000000}
};

localparam logic signed [12:0] bias [64] = '{
13'b1111111111101,  // -0.037350185215473175
13'b0000000010001,  // 0.27355897426605225
13'b1111111111000,  // -0.12378914654254913
13'b1111111111011,  // -0.064457006752491
13'b0000000000011,  // 0.05452875792980194
13'b0000000000111,  // 0.11671770364046097
13'b0000000001000,  // 0.13640816509723663
13'b0000000000100,  // 0.07482525706291199
13'b0000000000010,  // 0.04674031585454941
13'b1111111110011,  // -0.20146161317825317
13'b1111111111001,  // -0.09910125285387039
13'b0000000001001,  // 0.15104414522647858
13'b1111111111001,  // -0.10221704095602036
13'b1111111110110,  // -0.1461549550294876
13'b1111111111010,  // -0.08641516417264938
13'b0000000001010,  // 0.16613510251045227
13'b1111111111010,  // -0.0836295336484909
13'b1111111111100,  // -0.05756539851427078
13'b1111111111101,  // -0.03229188174009323
13'b1111111111110,  // -0.028388574719429016
13'b0000000001000,  // 0.1260243058204651
13'b1111111111101,  // -0.037064336240291595
13'b0000000001100,  // 0.19336333870887756
13'b0000000000001,  // 0.02124214917421341
13'b0000000011111,  // 0.4985624849796295
13'b0000000000001,  // 0.0158411655575037
13'b1111111111010,  // -0.08296407759189606
13'b0000000000111,  // 0.11056788265705109
13'b0000000000000,  // 0.01173810102045536
13'b1111111111001,  // -0.10843746364116669
13'b0000000010001,  // 0.27439257502555847
13'b0000000000101,  // 0.09199801832437515
13'b0000000010001,  // 0.27419957518577576
13'b0000000010001,  // 0.27063727378845215
13'b1111111110000,  // -0.24828937649726868
13'b0000000000101,  // 0.07818280160427094
13'b1111111111111,  // -0.005749030504375696
13'b0000000000110,  // 0.10850494354963303
13'b0000000001000,  // 0.13591453433036804
13'b1111111111000,  // -0.12088628858327866
13'b1111111111100,  // -0.05666546896100044
13'b0000000000101,  // 0.09311636537313461
13'b0000000000011,  // 0.05477767437696457
13'b0000000000001,  // 0.029585206881165504
13'b1111111101100,  // -0.31209176778793335
13'b1111111111010,  // -0.08465463668107986
13'b1111111110101,  // -0.16775836050510406
13'b0000000001001,  // 0.14762157201766968
13'b1111111110000,  // -0.23618532717227936
13'b0000000000100,  // 0.06535740196704865
13'b1111111110111,  // -0.12853026390075684
13'b1111111110111,  // -0.13802281022071838
13'b1111111110110,  // -0.15156887471675873
13'b0000000000101,  // 0.07979883998632431
13'b0000000001011,  // 0.18141601979732513
13'b1111111111100,  // -0.054039113223552704
13'b1111111111111,  // -0.010052933357656002
13'b0000000000100,  // 0.06611225008964539
13'b0000000000011,  // 0.05053366720676422
13'b0000000000001,  // 0.026860840618610382
13'b0000000000010,  // 0.03283466026186943
13'b0000000001001,  // 0.15558314323425293
13'b1111111101101,  // -0.2863388657569885
13'b1111111111010   // -0.08769102394580841
};
endpackage