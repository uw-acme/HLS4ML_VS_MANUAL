package reluDATA;

// For denseLatency
// RELU
localparam logic signed [16:0] weights[0:319] = '{
17'b00000000011110000,
17'b11111111101000000,
17'b00000000000100001,
17'b11111111111001111,
17'b11111111010000001,
17'b00000001010010110,
17'b00000000000110011,
17'b00000000101000000,
17'b00000000101011010,
17'b11111111110000110,
17'b11111111110010101,
17'b11111111111111100,
17'b00000000001000011,
17'b00000000011001000,
17'b00000000000011011,
17'b00000000100001001,
17'b11111111111011000,
17'b11111111110010001,
17'b11111111011000010,
17'b00000000010001001,
17'b00000000101000010,
17'b00000000000111110,
17'b11111110110010001,
17'b00000000011011010,
17'b00000000000011111,
17'b00000000001110010,
17'b00000000101011001,
17'b11111110111111011,
17'b00000000111010111,
17'b00000000010010100,
17'b00000001001011100,
17'b11111111101110010,
17'b00000000111110101,
17'b00000001110110111,
17'b11111111110110100,
17'b00000000001101101,
17'b00000000010110011,
17'b00000000000101110,
17'b11111111111110100,
17'b00000000100010001,
17'b00000000011011110,
17'b11111111111001001,
17'b00000001000010101,
17'b00000001011110111,
17'b00000000011010001,
17'b00000000011000010,
17'b00000001011000111,
17'b11111111111010000,
17'b11111111111000010,
17'b11111111010011111,
17'b11111111100001011,
17'b00000000011001011,
17'b11111111101011101,
17'b00000000011111001,
17'b00000001000111101,
17'b11111111111000110,
17'b11111111011001100,
17'b00000000010001111,
17'b00000001111011010,
17'b11111111111111100,
17'b00000000000010010,
17'b11111110110100000,
17'b11111111001001110,
17'b00000000011001110,
17'b11111101010110100,
17'b11111110100011100,
17'b11111101101111110,
17'b00000000011001001,
17'b11111111001010111,
17'b00000001100001110,
17'b11111111010110001,
17'b11111111010011000,
17'b00000000000011001,
17'b11111101001100101,
17'b11111111001011111,
17'b11111110011100010,
17'b11111111101000011,
17'b11111111010010111,
17'b11111111001101001,
17'b00000000100110011,
17'b00000001001011111,
17'b00000000011100001,
17'b11111110001100010,
17'b00000000110011101,
17'b00000001010011100,
17'b00000000100110111,
17'b11111111100010100,
17'b00000001010110111,
17'b11111110101000001,
17'b00000001000100110,
17'b00000000111001001,
17'b00000000110011110,
17'b11111111101100011,
17'b11111111111000101,
17'b11111111101100010,
17'b11111111111111011,
17'b11111110000100011,
17'b11111110100010101,
17'b00000000001001011,
17'b11111111101111110,
17'b11111111101010001,
17'b00000001011110001,
17'b00000000111101010,
17'b11111111110011000,
17'b00000000010100110,
17'b11111111011111011,
17'b00000000000010110,
17'b11111110111100111,
17'b11111110011101110,
17'b11111111101110000,
17'b00000000110000001,
17'b00000000111110001,
17'b00000000111010101,
17'b11111110110011000,
17'b11111110111110000,
17'b11111111011000111,
17'b00000000100110001,
17'b11111110110111100,
17'b00000000010010000,
17'b11111111011101111,
17'b11111111011000001,
17'b00000000101110000,
17'b11111111111100100,
17'b00000001010111000,
17'b11111111111010001,
17'b11111110110110111,
17'b11111111101100010,
17'b00000000100110001,
17'b00000000000110010,
17'b00000000101000010,
17'b11111111100100000,
17'b00000001010110100,
17'b00000000011101000,
17'b11111111010001000,
17'b00000000010110001,
17'b00000000101100000,
17'b00000001010101100,
17'b11111111010000011,
17'b11111111111110101,
17'b11111111011010101,
17'b00000000101111000,
17'b00000000100100110,
17'b00000000010001011,
17'b11111111010010100,
17'b11111111011111101,
17'b00000000011101111,
17'b11111110100011011,
17'b00000000010111111,
17'b00000000011010111,
17'b00000000010111000,
17'b11111111010100111,
17'b11111111101000010,
17'b00000000001110011,
17'b11111111001111011,
17'b11111111100010010,
17'b11111111110101100,
17'b11111111000001101,
17'b00000000101101001,
17'b00000000111111111,
17'b11111111100110000,
17'b00000000000011000,
17'b11111111010011111,
17'b11111111001011000,
17'b00000001010010100,
17'b11111110101110101,
17'b00000000000000101,
17'b11111111101110100,
17'b11111111101000101,
17'b00000000010001001,
17'b00000000010010100,
17'b00000000010001000,
17'b00000000100110001,
17'b11111111111011110,
17'b11111111101000110,
17'b11111111011000110,
17'b11111111011011101,
17'b00000001000111101,
17'b00000001000001111,
17'b11111111011001111,
17'b00000001001000100,
17'b00000000010000000,
17'b00000000001011111,
17'b00000000101011111,
17'b00000000110101110,
17'b11111111100010110,
17'b00000000101110110,
17'b11111111101111001,
17'b11111111100100001,
17'b11111111011101101,
17'b11111111010110111,
17'b11111111000000101,
17'b00000000010010100,
17'b11111111111010101,
17'b00000001001110000,
17'b11111111010100001,
17'b11111111101011010,
17'b00000000100111011,
17'b11111111111011100,
17'b00000000111110111,
17'b00000000011100100,
17'b00000000100000011,
17'b00000000110011101,
17'b00000001001101011,
17'b00000001001011010,
17'b00000000011101011,
17'b11111111110101101,
17'b00000000100100010,
17'b11111111001100000,
17'b11111110110010011,
17'b11111110100101110,
17'b00000001001010100,
17'b00000001001111001,
17'b11111111001101100,
17'b00000000010100010,
17'b11111111111101111,
17'b00000000010100101,
17'b00000000011111011,
17'b00000001001111110,
17'b11111111101001011,
17'b00000000000001010,
17'b00000001100001000,
17'b11111111000011111,
17'b11111111101010101,
17'b11111110000000001,
17'b00000001001000000,
17'b00000000100111110,
17'b00000001011100111,
17'b11111111100111001,
17'b00000000011100010,
17'b11111111001000001,
17'b11111111100000110,
17'b11111111100000000,
17'b11111111100100110,
17'b00000000001111000,
17'b00000001000110000,
17'b00000000010111001,
17'b11111111111001001,
17'b00000000001011011,
17'b11111111111111110,
17'b00000000010110110,
17'b11111111011000011,
17'b00000000000001010,
17'b00000000001111100,
17'b00000001001110000,
17'b11111111001011100,
17'b00000000110111010,
17'b00000000010111000,
17'b11111111001111001,
17'b00000000100101011,
17'b11111111001110010,
17'b00000000010101010,
17'b11111111000100010,
17'b00000001001111110,
17'b11111111011100101,
17'b11111111011010111,
17'b11111111000010000,
17'b00000010000000100,
17'b00000000101100011,
17'b00000000010100001,
17'b00000000011000100,
17'b11111111110111000,
17'b11111111110000101,
17'b00000001001100000,
17'b00000001000110010,
17'b11111111111101010,
17'b00000000110010011,
17'b00000001000011110,
17'b11111101011011100,
17'b00000010010010101,
17'b11111100100000111,
17'b11111110100101101,
17'b11111111101000100,
17'b11111111111010011,
17'b00000001010101111,
17'b00000000001000111,
17'b11111111011101100,
17'b00000000100010101,
17'b00000001101110110,
17'b00000000011111000,
17'b11111111110000001,
17'b00000000101000100,
17'b11111111000100111,
17'b11111110110010100,
17'b11111110110110111,
17'b00000000101011000,
17'b00000001110111011,
17'b00000000111010111,
17'b11111101110000000,
17'b11111111001010010,
17'b11111110111101110,
17'b11111111111011100,
17'b00000001100000000,
17'b00000000100110011,
17'b00000000011110101,
17'b11111111000101001,
17'b11111110000101011,
17'b00000001011000101,
17'b11111110110001111,
17'b11111111000110100,
17'b11111101110111001,
17'b11111111101111010,
17'b00000000011000011,
17'b11111111010110110,
17'b11111111010010111,
17'b00000001000010101,
17'b00000001000100101,
17'b11111111110011010,
17'b11111111001111000,
17'b00000000111010100,
17'b00000001101100001,
17'b00000000101100100,
17'b00000001110001110,
17'b11111111000011011,
17'b00000001100111101,
17'b00000000000110001,
17'b00000000001011101,
17'b11111111111100110,
17'b00000000011011001,
17'b11111111101011011,
17'b00000000000101010
};

localparam logic signed [16:0] bias[0:31] = '{
17'b00000001101011110,
17'b00000001100101001,
17'b00000001010011000,
17'b00000000001001000,
17'b00000000110100010,
17'b00000000000000000,
17'b11111111001111010,
17'b00000000111100101,
17'b00000000000000100,
17'b00000001110011101,
17'b00000000110100111,
17'b00000000100101010,
17'b00000000010111111,
17'b00000001100011001,
17'b00000001111101100,
17'b11111111111011110,
17'b00000000010001011,
17'b11111110111111000,
17'b00000000100011110,
17'b11111111101011000,
17'b00000000001110101,
17'b00000000111011001,
17'b00000000000110111,
17'b11111111011100010,
17'b00000001101110011,
17'b11111111111111011,
17'b00000000110111011,
17'b00000000001101111,
17'b00000000111001100,
17'b00000000100010100,
17'b00000001000000111,
17'b11111111111100111
};
endpackage
