// Width: 18
// NFRAC: 9
package dense_2_18_9;

localparam logic signed [17:0] weights [64][32] = '{ 
{18'b000000000010001001, 18'b000000000000000100, 18'b111111111110011110, 18'b111111111111110101, 18'b000000000010000101, 18'b000000000000000000, 18'b111111111110110110, 18'b111111111111111111, 18'b111111111101110011, 18'b000000000000101000, 18'b000000000000000000, 18'b111111111111111101, 18'b111111111111111111, 18'b111111111110011001, 18'b111111111111100110, 18'b111111111101111001, 18'b000000000000000000, 18'b111111111111111001, 18'b111111111110011110, 18'b111111111110101110, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111111111011, 18'b111111111111111110, 18'b000000000000000000, 18'b000000000000110011, 18'b000000000011000101, 18'b000000000001011001, 18'b111111111111111111, 18'b000000000000011001, 18'b111111111100101110, 18'b000000000000000000}, 
{18'b111111111111001100, 18'b111111111110110000, 18'b111111111110111001, 18'b111111111111100011, 18'b111111111111111101, 18'b000000000000010110, 18'b111111111110001101, 18'b000000000000000010, 18'b000000000000000010, 18'b111111111111011111, 18'b000000000001001111, 18'b111111111111101001, 18'b111111111111100001, 18'b111111111110010000, 18'b000000000000000011, 18'b111111111111100111, 18'b000000000000000110, 18'b111111111110011100, 18'b000000000001010111, 18'b000000000001110101, 18'b111111111111101111, 18'b111111111111111101, 18'b111111111111111111, 18'b000000000000001100, 18'b111111111111011011, 18'b000000000010001100, 18'b000000000001111110, 18'b000000000000000100, 18'b000000000000001110, 18'b111111111100000110, 18'b000000000000000011, 18'b000000000000000000}, 
{18'b000000000000100101, 18'b111111111111000101, 18'b111111111110111101, 18'b111111111111101010, 18'b111111111111011000, 18'b111111111111010100, 18'b111111111110100001, 18'b000000000000000010, 18'b111111111110111010, 18'b000000000000000100, 18'b000000000000000001, 18'b111111111111010110, 18'b000000000000101110, 18'b111111111111011110, 18'b111111111111111111, 18'b111111111111101101, 18'b000000000000000010, 18'b000000000000110000, 18'b000000000000011110, 18'b000000000001110101, 18'b000000000000010101, 18'b111111111111010100, 18'b000000000000000000, 18'b000000000000010001, 18'b111111111111110110, 18'b000000000001101011, 18'b000000000001001100, 18'b000000000000110001, 18'b111111111111111111, 18'b111111111110110010, 18'b111111111111111001, 18'b000000000000110010}, 
{18'b000000000001000110, 18'b000000000000001001, 18'b000000000000011011, 18'b111111111111111011, 18'b111111111011111011, 18'b000000000000000000, 18'b000000000000000000, 18'b000000000001110011, 18'b000000000001111100, 18'b111111111111111001, 18'b111111111111111111, 18'b000000000000000000, 18'b000000000000000000, 18'b000000000000000010, 18'b111111111111110110, 18'b000000000001101101, 18'b000000000000000000, 18'b111111111111110011, 18'b111111111111111111, 18'b111111111110100101, 18'b111111111111100000, 18'b000000000000011001, 18'b111111111111011111, 18'b111111111111111111, 18'b000000000000000001, 18'b111111111111100110, 18'b000000000000100101, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111110010001, 18'b000000000010011110}, 
{18'b111111111010100010, 18'b111111111111110011, 18'b111111111111111101, 18'b000000000000000010, 18'b111111111111110010, 18'b000000000000000011, 18'b111111111111100110, 18'b111111111110110011, 18'b000000000000011011, 18'b111111111111110101, 18'b111111111111111001, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000001101011, 18'b000000000000000000, 18'b000000000010101000, 18'b111111111111111111, 18'b000000000001101111, 18'b111111111100110011, 18'b000000000000000000, 18'b111111111111000110, 18'b000000000001010110, 18'b000000000010000100, 18'b000000000000000000, 18'b000000000000010111, 18'b000000000001010011, 18'b000000000001111010, 18'b000000000000001000, 18'b111111111111111101, 18'b111111111111111111, 18'b111111111111111000, 18'b000000000001110011}, 
{18'b000000000000011101, 18'b111111111111111111, 18'b000000000001001100, 18'b111111111010110011, 18'b111111110100111110, 18'b111111111101001100, 18'b000000000010110101, 18'b111111111011000001, 18'b111111111111111111, 18'b111111111010100101, 18'b111111111011111111, 18'b111111111101010001, 18'b000000000010110100, 18'b111111111111111111, 18'b111111111111111000, 18'b000000000000000000, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111110111100, 18'b111111111111111111, 18'b111111111100000101, 18'b000000000000000000, 18'b000000000001011111, 18'b111111111111111111, 18'b000000000000001011, 18'b000000000010001001, 18'b000000000000011010, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000001101001, 18'b111111111111101110, 18'b000000000001100110}, 
{18'b111111111111101101, 18'b111111111110101111, 18'b111111111110000100, 18'b111111111111100111, 18'b111111111101101100, 18'b000000000000100001, 18'b111111111110100011, 18'b111111111110110111, 18'b111111111100101011, 18'b000000000000011000, 18'b111111111111111101, 18'b111111111110101110, 18'b000000000000111100, 18'b111111111111111010, 18'b111111111111101010, 18'b111111111011100100, 18'b111111111111111111, 18'b000000000000101011, 18'b000000000001100010, 18'b111111111110101100, 18'b111111111110110011, 18'b111111111111011111, 18'b111111111111111111, 18'b000000000000001110, 18'b111111111111101000, 18'b111111111010110100, 18'b111111111101111000, 18'b111111111111101000, 18'b000000000000000010, 18'b111111111111110101, 18'b000000000000001111, 18'b111111111111111111}, 
{18'b111111111110110001, 18'b111111111111010001, 18'b111111111111010111, 18'b111111111110000110, 18'b111111111111000100, 18'b111111111111111111, 18'b000000000000110101, 18'b111111111111010111, 18'b000000000001100110, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111111111111, 18'b000000000001110000, 18'b000000000000000000, 18'b111111111111111111, 18'b111111111111011011, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111111111111, 18'b000000000000010110, 18'b111111111110100011, 18'b000000000000000111, 18'b111111111111111111, 18'b111111111111011011, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111111111111}, 
{18'b111111111100001011, 18'b111111111111100010, 18'b111111111100111101, 18'b000000000000111110, 18'b000000000011111001, 18'b111111111111111111, 18'b111111111111110001, 18'b000000000001111010, 18'b111111111100011111, 18'b111111111111101000, 18'b000000000000000000, 18'b111111111110011000, 18'b111111111111111111, 18'b000000000000100110, 18'b111111111110011110, 18'b000000000110000010, 18'b111111111111111011, 18'b000000000000010111, 18'b000000000001101010, 18'b000000000001111101, 18'b000000000000000000, 18'b111111111101010100, 18'b000000000000000000, 18'b000000000011010010, 18'b111111111110100011, 18'b000000000101100101, 18'b111111111110110011, 18'b111111111110010111, 18'b111111111100001110, 18'b111111111100010010, 18'b000000000000000000, 18'b000000000000011011}, 
{18'b000000000000000000, 18'b111111111111111000, 18'b111111111111011010, 18'b000000000000000000, 18'b000000000010011101, 18'b111111111111110101, 18'b111111111111011111, 18'b000000000000101111, 18'b000000000000110011, 18'b000000000000000001, 18'b111111111111111011, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111111000101, 18'b111111111111111111, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111111111101, 18'b000000000000000001, 18'b000000000000101011, 18'b000000000000001001, 18'b111111111111111111, 18'b000000000000000000, 18'b000000000000000011, 18'b000000000000010011, 18'b111111111110111100, 18'b000000000000100010, 18'b000000000001111111, 18'b111111111111111111, 18'b000000000000000011, 18'b000000000000011001, 18'b000000000000100011}, 
{18'b000000000000110001, 18'b000000000000000000, 18'b111111111111001011, 18'b111111111101111111, 18'b111111111001101001, 18'b000000000001000100, 18'b000000000000000000, 18'b111111111001011000, 18'b000000000000010010, 18'b111111111111111111, 18'b000000000000000001, 18'b111111111111111111, 18'b000000000000000101, 18'b000000000000000000, 18'b111111111111110110, 18'b111111111100111100, 18'b111111111111111111, 18'b000000000001110000, 18'b000000000001000000, 18'b000000000001100001, 18'b111111111100011110, 18'b111111111101001001, 18'b000000000000111101, 18'b111111111111101110, 18'b111111111111101000, 18'b000000000010110111, 18'b111111111111001110, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000001101100, 18'b111111111111111111, 18'b000000000000000011}, 
{18'b111111111110011010, 18'b111111111100000011, 18'b000000000000000000, 18'b111111111111111110, 18'b000000000010101010, 18'b111111111101110110, 18'b111111111110001110, 18'b000000000000111011, 18'b111111111111111111, 18'b000000000001001100, 18'b000000000000100101, 18'b111111111111011001, 18'b000000000000000000, 18'b000000000000000111, 18'b111111111111110101, 18'b111111111101111110, 18'b000000000001011001, 18'b000000000000001110, 18'b000000000010011000, 18'b000000000000101100, 18'b000000000000000000, 18'b111111111111101100, 18'b000000000001000000, 18'b111111111111010011, 18'b111111111101100010, 18'b111111111111111100, 18'b000000000001011110, 18'b111111111111111111, 18'b000000000000000100, 18'b111111111111001111, 18'b000000000001000110, 18'b000000000010001101}, 
{18'b000000000000000111, 18'b000000000000000000, 18'b000000000001110000, 18'b000000000000000100, 18'b111111111111101011, 18'b000000000001011100, 18'b000000000000101111, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111110111000, 18'b111111111111100100, 18'b111111111110101010, 18'b111111111111111111, 18'b000000000000011001, 18'b111111111111011100, 18'b000000000110101111, 18'b000000000000000000, 18'b111111111111001111, 18'b111111111110011111, 18'b111111111111111001, 18'b000000000001100101, 18'b000000000001000001, 18'b000000000000000000, 18'b111111111111111110, 18'b000000000001110000, 18'b000000000010001001, 18'b000000000011111101, 18'b000000000000000101, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111111111001, 18'b111111111111011011}, 
{18'b111111111110110000, 18'b000000000000011000, 18'b000000000000010100, 18'b111111111110000001, 18'b111111111101110110, 18'b000000000011110000, 18'b000000000000011001, 18'b000000000000000000, 18'b111111111110101101, 18'b111111111111010010, 18'b000000000001000010, 18'b000000000000100100, 18'b000000000000000000, 18'b111111111111010111, 18'b000000000010010010, 18'b111111111111111111, 18'b111111111111111001, 18'b000000000000000000, 18'b000000000000000110, 18'b111111111111101000, 18'b000000000000101000, 18'b000000000000001000, 18'b000000000000111010, 18'b111111111111111111, 18'b000000000000000001, 18'b000000000101010000, 18'b111111111111100011, 18'b111111111111110100, 18'b111111111111111111, 18'b111111111111001000, 18'b111111111111101011, 18'b000000000001011010}, 
{18'b000000000000011110, 18'b000000000000100101, 18'b000000000010100111, 18'b111111111111101011, 18'b000000000000110011, 18'b000000000010110011, 18'b000000000000000000, 18'b111111111111110000, 18'b000000000000111100, 18'b111111111111000101, 18'b111111111111111111, 18'b111111111111000010, 18'b000000000000000000, 18'b000000000011001001, 18'b111111111111110110, 18'b000000000000000000, 18'b000000000001111000, 18'b000000000000000000, 18'b000000000000000001, 18'b111111111101011111, 18'b111111111110000010, 18'b111111111111101101, 18'b111111111111111111, 18'b111111111110110101, 18'b111111111111101101, 18'b111111111111010101, 18'b111111111110011011, 18'b111111111110010011, 18'b000000000000001111, 18'b000000000000111001, 18'b111111111100110100, 18'b000000000000000001}, 
{18'b111111111101100111, 18'b000000000000000000, 18'b111111111111111000, 18'b111111111111100110, 18'b111111111111111111, 18'b000000000001000100, 18'b111111111111011000, 18'b000000000010001010, 18'b111111111101000110, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111111111111, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111111111110, 18'b111111111111010001, 18'b000000000000101000, 18'b000000000001011101, 18'b111111111111111011, 18'b111111111101111111, 18'b111111111111100001, 18'b000000000000111001, 18'b000000000000100000, 18'b000000000000000000, 18'b000000000000000001, 18'b000000000000101001, 18'b111111111110000101, 18'b000000000000000000, 18'b111111111111111111, 18'b000000000000000001, 18'b000000000000000000, 18'b111111111110111111}, 
{18'b111111111101010011, 18'b111111111111111101, 18'b111111111111111110, 18'b111111111111110111, 18'b111111111111111101, 18'b000000000000110110, 18'b000000000000000011, 18'b000000000000010001, 18'b000000000000010011, 18'b000000000000100000, 18'b000000000000101000, 18'b000000000001010010, 18'b000000000000001101, 18'b111111111111001110, 18'b000000000000000000, 18'b000000000011000011, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111111111110, 18'b000000000000111000, 18'b000000000001001000, 18'b000000000000001111, 18'b000000000000010101, 18'b111111111111110000, 18'b111111111111101111, 18'b000000000000001101, 18'b111111111111011101, 18'b111111111110111111, 18'b000000000001101011, 18'b111111111111110000, 18'b000000000000010000, 18'b111111111110011111}, 
{18'b000000000000000000, 18'b111111111111111111, 18'b000000000000010011, 18'b000000000000000000, 18'b000000000111010000, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111111111111, 18'b000000000000111000, 18'b111111111111011001, 18'b000000000000000000, 18'b000000000000000000, 18'b000000000000000000, 18'b000000000001000010, 18'b000000000000000000, 18'b111111111110110101, 18'b111111111111111111, 18'b111111111111011101, 18'b000000000010100111, 18'b000000000000000000, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111111111111, 18'b000000000000000000, 18'b000000000000100010, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000000000000, 18'b000000000000010101}, 
{18'b111111111111111110, 18'b000000000000001110, 18'b111111111111111111, 18'b000000000000011000, 18'b111111111111101001, 18'b111111111111000010, 18'b111111111111100000, 18'b000000000010001110, 18'b000000000000000000, 18'b000000000000110001, 18'b111111111111111010, 18'b000000000000100001, 18'b111111111111101111, 18'b111111111110101111, 18'b111111111110011110, 18'b000000000000000110, 18'b111111111111111111, 18'b111111111111101110, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111111111111, 18'b000000000000100110, 18'b000000000000010010, 18'b111111111110111111, 18'b000000000000111001, 18'b111111111110101011, 18'b000000000000000001, 18'b000000000000000000, 18'b111111111110101010, 18'b000000000000000000, 18'b000000000000010111, 18'b111111111111110000}, 
{18'b111111111111111010, 18'b111111111111001101, 18'b000000000000000000, 18'b111111111111100001, 18'b000000000001101110, 18'b111111111111111111, 18'b111111111111110101, 18'b000000000000110110, 18'b111111111100110111, 18'b000000000000000000, 18'b111111111111101100, 18'b111111111111111110, 18'b000000000010110011, 18'b000000000001110101, 18'b111111111111001101, 18'b111111111111110101, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111111111111, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111110111010, 18'b111111111111000011, 18'b000000000001000011, 18'b000000000000000000, 18'b111111111110111001, 18'b000000000000001100, 18'b111111111111010110, 18'b111111111111101110, 18'b000000000001000101, 18'b000000000000000000, 18'b111111111110000001}, 
{18'b000000000101000100, 18'b000000000010101111, 18'b111111111110000000, 18'b000000000000000001, 18'b111111111101001110, 18'b000000000000000000, 18'b000000000001110010, 18'b000000000000001111, 18'b000000000001110010, 18'b111111111111111111, 18'b111111111110110000, 18'b111111111111010111, 18'b000000000001001000, 18'b000000000000001110, 18'b111111111111001101, 18'b000000000001000011, 18'b000000000100010010, 18'b111111111110111101, 18'b111111111101101000, 18'b000000000000000000, 18'b111111111111110001, 18'b111111111110100101, 18'b111111111111111001, 18'b111111111111111111, 18'b000000000000101100, 18'b111111111101000111, 18'b000000000000101101, 18'b111111111111111111, 18'b000000000000000000, 18'b000000000000110111, 18'b111111111111110001, 18'b000000000000011110}, 
{18'b111111111111010000, 18'b111111111110011101, 18'b111111111111101101, 18'b111111111110101010, 18'b111111111111110111, 18'b000000000000011001, 18'b000000000000000000, 18'b111111111111111010, 18'b000000000000010011, 18'b111111111111111110, 18'b000000000000000000, 18'b111111111110010000, 18'b000000000000110100, 18'b000000000000101001, 18'b111111111111001011, 18'b000000000011100011, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111111111101, 18'b000000000000000000, 18'b000000000010100001, 18'b111111111100001111, 18'b111111111111001000, 18'b111111111111100011, 18'b111111111111110110, 18'b000000000001100100, 18'b111111111111100101, 18'b000000000000001001, 18'b000000000011110111, 18'b111111111011111001, 18'b111111111101000100, 18'b000000000000001011}, 
{18'b000000000000001000, 18'b111111111111100001, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111010001111, 18'b111111111011001001, 18'b000000000000000000, 18'b111111111111111111, 18'b111111111101111000, 18'b000000000000001100, 18'b000000000000000000, 18'b111111111111110001, 18'b000000000000000000, 18'b111111111111100010, 18'b111111111111100101, 18'b111111111111011100, 18'b111111111110110100, 18'b000000000010010000, 18'b000000000000000000, 18'b000000000000010111, 18'b111111111111111111, 18'b111111111111011011, 18'b000000000000000000, 18'b111111111111010011, 18'b000000000001110000, 18'b111111111011000001, 18'b000000000001110000, 18'b111111111111111111, 18'b111111111111111101, 18'b000000000001100110, 18'b111111111111111111, 18'b000000000001111000}, 
{18'b111111111111111111, 18'b000000000000000010, 18'b111111111111101001, 18'b000000000000100110, 18'b000000000000011100, 18'b111111111101010000, 18'b000000000000000000, 18'b000000000000100000, 18'b000000000100101000, 18'b111111111111111011, 18'b000000000000000000, 18'b000000000000011100, 18'b000000000010110111, 18'b111111111111101111, 18'b000000000000000111, 18'b000000000000110011, 18'b111111111111111111, 18'b000000000000001110, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111101110011, 18'b000000000000010011, 18'b000000000000100011, 18'b000000000000001011, 18'b111111111111111111, 18'b000000000001101111, 18'b000000000000000010, 18'b000000000001000000, 18'b111111111100101010, 18'b000000000000110100, 18'b000000000011001010, 18'b000000000000000010}, 
{18'b111111111101001100, 18'b000000000001101100, 18'b111111111101111010, 18'b000000000000111110, 18'b111111111111001010, 18'b000000000000000000, 18'b000000000011111110, 18'b111111111110001000, 18'b111111111101101010, 18'b000000000001010111, 18'b111111111110001101, 18'b111111111111110011, 18'b111111111111111111, 18'b000000000010110000, 18'b111111111111111111, 18'b111111111101100101, 18'b111111111111111111, 18'b000000000011100001, 18'b111111111100001110, 18'b111111111111110011, 18'b000000000010100010, 18'b111111111101000110, 18'b000000000000011011, 18'b111111111111111000, 18'b000000000010001010, 18'b111111111011111011, 18'b111111111101000110, 18'b111111111110011011, 18'b111111111111111111, 18'b000000000000110101, 18'b000000000000001100, 18'b000000000001011011}, 
{18'b111111111111010001, 18'b000000000000011010, 18'b111111111111111111, 18'b000000000001001100, 18'b111111111111101100, 18'b000000000001110100, 18'b000000000000000001, 18'b111111111111111010, 18'b111111111111111110, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000100001010, 18'b000000000000000110, 18'b000000000001100000, 18'b000000000000000000, 18'b111111111110010011, 18'b111111111111011000, 18'b111111111111111111, 18'b111111111111110111, 18'b000000000000010101, 18'b111111111111111111, 18'b111111111110100001, 18'b111111111111111111, 18'b000000000010010111, 18'b000000000010011110, 18'b111111111111111111, 18'b111111111111110111, 18'b000000000000000000, 18'b111111111111111111, 18'b111111111111001110}, 
{18'b111111111111010110, 18'b000000000000000000, 18'b000000000010001011, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111111000101, 18'b000000000000000000, 18'b111111111001000101, 18'b000000000001101110, 18'b000000000000000111, 18'b000000000000001101, 18'b111111111101000111, 18'b000000000000000001, 18'b111111111110111001, 18'b111111111111101111, 18'b000000000000000000, 18'b000000000000001010, 18'b000000000000000000, 18'b000000000000111001, 18'b000000000000000000, 18'b111111111111111011, 18'b000000000010101000, 18'b000000000011000000, 18'b111111111110001110, 18'b111111111110110111, 18'b000000000001111111, 18'b111111111101100011, 18'b000000000000001111, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000001011110}, 
{18'b111111111111000101, 18'b111111111111111111, 18'b111111111110000101, 18'b111111111110011000, 18'b111111111111111000, 18'b111111111110111010, 18'b000000000000000000, 18'b000000000000101110, 18'b111111111110000101, 18'b111111111111010101, 18'b111111111111100110, 18'b000000000000000000, 18'b000000000000001110, 18'b111111111111111010, 18'b111111111111100000, 18'b000000000000110000, 18'b000000000001110010, 18'b000000000001000011, 18'b111111111110111101, 18'b000000000000011000, 18'b111111111111111001, 18'b111111111111110001, 18'b000000000000001011, 18'b000000000000001000, 18'b111111111111011100, 18'b000000000000101101, 18'b111111111111010001, 18'b000000000000011110, 18'b111111111111111111, 18'b111111111101101000, 18'b111111111111110010, 18'b000000000001110011}, 
{18'b111111111111110010, 18'b111111111111010101, 18'b000000000000100111, 18'b000000000010000001, 18'b000000000000101011, 18'b000000000000101010, 18'b000000000000010111, 18'b111111111110011000, 18'b111111111110010110, 18'b000000000000100011, 18'b000000000000000110, 18'b000000000000010110, 18'b000000000000001011, 18'b000000000000000010, 18'b000000000001101001, 18'b000000000000000011, 18'b111111111111100100, 18'b000000000000110100, 18'b111111111111110000, 18'b111111111111101101, 18'b000000000000111000, 18'b111111111111000000, 18'b111111111111110010, 18'b000000000001000001, 18'b000000000000001011, 18'b111111111111001001, 18'b111111111110011010, 18'b111111111111111001, 18'b111111111101110001, 18'b000000000000011110, 18'b000000000000110100, 18'b000000000000000000}, 
{18'b111111111111111001, 18'b111111111111110101, 18'b111111111111111001, 18'b111111111111101110, 18'b111111111110111100, 18'b111111111110111000, 18'b000000000000100000, 18'b000000000000000100, 18'b111111111110100010, 18'b000000000001010101, 18'b111111111111110101, 18'b111111111111111111, 18'b111111111111000111, 18'b000000000000000010, 18'b000000000000001111, 18'b111111111111100101, 18'b111111111111110111, 18'b111111111111101010, 18'b111111111111010110, 18'b000000000000000000, 18'b111111111110111000, 18'b000000000000110100, 18'b111111111110010011, 18'b000000000000000010, 18'b000000000000010101, 18'b000000000000111111, 18'b000000000000001101, 18'b000000000000000011, 18'b000000000010010101, 18'b000000000000011010, 18'b000000000000000000, 18'b000000000000101010}, 
{18'b111111111111110110, 18'b000000000010000001, 18'b111111111111111111, 18'b111111111111101111, 18'b111111111110010010, 18'b111111111111011001, 18'b000000000011010010, 18'b111111111010011111, 18'b111111111101001101, 18'b111111111110011001, 18'b111111111110001111, 18'b111111111101111110, 18'b111111111111111111, 18'b000000000011110111, 18'b111111111111110010, 18'b000000000000000000, 18'b111111111110010011, 18'b000000000011100100, 18'b111111111100101100, 18'b000000000000000000, 18'b111111111111111111, 18'b111111111101010011, 18'b000000000000000000, 18'b111111111111111111, 18'b000000000000011100, 18'b111111111111100010, 18'b111111111110110100, 18'b111111111111111111, 18'b000000000001011001, 18'b000000000000000001, 18'b111111111111010110, 18'b000000000000000000}, 
{18'b000000000010111100, 18'b111111111111000110, 18'b000000000001000011, 18'b111111111111101111, 18'b000000000000100111, 18'b111111111111111110, 18'b111111111111111110, 18'b111111111111010000, 18'b000000000000000000, 18'b000000000000101111, 18'b111111111111111111, 18'b111111111111100001, 18'b111111111111111111, 18'b000000000001110101, 18'b000000000000001001, 18'b000000000000010100, 18'b000000000000001100, 18'b111111111111110011, 18'b000000000000001010, 18'b000000000000000000, 18'b111111111111111011, 18'b111111111111111111, 18'b111111111101100011, 18'b111111111111111111, 18'b000000000000011101, 18'b111111111111000100, 18'b111111111110111010, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000100011101, 18'b111111111101101101, 18'b111111111111000100}, 
{18'b111111111111101001, 18'b111111111111001011, 18'b111111111111011110, 18'b000000000000010010, 18'b000000000001000111, 18'b111111111110111101, 18'b111111111111111111, 18'b111111111110001111, 18'b000000000000011111, 18'b000000000001000101, 18'b111111111110010010, 18'b111111111101111110, 18'b000000000000001100, 18'b111111111010100010, 18'b111111111111011001, 18'b111111111111000000, 18'b111111111110011010, 18'b111111111111111111, 18'b000000000001000100, 18'b000000000000000000, 18'b111111111111101000, 18'b111111111111101001, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111111100001, 18'b111111111001111101, 18'b111111111011100011, 18'b111111111101110100, 18'b000000000000011100, 18'b000000000001101001, 18'b111111111111111111, 18'b000000000001111011}, 
{18'b111111111111010000, 18'b111111111110010010, 18'b000000000001010011, 18'b000000000000100110, 18'b000000000000010110, 18'b111111111111010000, 18'b111111111111101111, 18'b000000000000110010, 18'b000000000100010011, 18'b111111111110101000, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000000111100, 18'b111111111111100011, 18'b111111111111110110, 18'b111111111111110111, 18'b111111111111001100, 18'b111111111111111111, 18'b000000000000000000, 18'b000000000001110100, 18'b111111111110111011, 18'b111111111111111110, 18'b000000000001000001, 18'b111111111111111010, 18'b000000000000000000, 18'b000000000100001101, 18'b000000000010100110, 18'b000000000000000001, 18'b000000000000000000, 18'b111111111100101000, 18'b111111111111011101, 18'b111111111111111111}, 
{18'b000000000000000111, 18'b000000000000011000, 18'b111111111111111000, 18'b000000000000000000, 18'b000000000001110110, 18'b111111111100001000, 18'b000000000000000000, 18'b111111111111001111, 18'b000000000001011111, 18'b000000000000000000, 18'b111111111111110110, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111111111111, 18'b000000000000000010, 18'b111111111111001000, 18'b000000000010000100, 18'b111111111111111101, 18'b111111111111111000, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111111111100, 18'b000000000000000000, 18'b111111111111111111, 18'b000000000000000110, 18'b111111111101011101, 18'b000000000000011010, 18'b000000000001011101, 18'b111111111111111110, 18'b000000000000110000, 18'b111111111111111111, 18'b000000000000100110}, 
{18'b111111111110011000, 18'b000000000000000100, 18'b111111111100001001, 18'b000000000000000011, 18'b111111111111100110, 18'b111111111111101011, 18'b111111111111111111, 18'b111111111111010001, 18'b111111111111101101, 18'b111111111111011110, 18'b000000000000011000, 18'b000000000000001101, 18'b111111111110100101, 18'b000000000000000000, 18'b111111111111111111, 18'b111111111111111011, 18'b000000000000100100, 18'b111111111111110101, 18'b111111111111110001, 18'b111111111111110001, 18'b111111111111111111, 18'b000000000010001010, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111111111011, 18'b000000000010100010, 18'b000000000001100000, 18'b000000000000010001, 18'b111111111111001110, 18'b111111111111111010, 18'b000000000000100001, 18'b000000000000011101}, 
{18'b000000000000010001, 18'b000000000000010100, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111100010000, 18'b000000000000010110, 18'b000000000000001100, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111110101001, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111110101101, 18'b000000000000000000, 18'b000000000000000000, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111101001001, 18'b000000000000000100, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000000000000, 18'b000000000001000010, 18'b111111111111111111, 18'b000000000000000000, 18'b000000000011101001, 18'b000000000010101110, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111110001000, 18'b000000000000000000, 18'b111111111111111111}, 
{18'b000000000000100110, 18'b000000000000011011, 18'b000000000010000001, 18'b111111111110000000, 18'b000000000001000011, 18'b000000000000111100, 18'b000000000000000011, 18'b000000000001100010, 18'b000000000000000110, 18'b111111111111111001, 18'b000000000000010011, 18'b000000000000000010, 18'b111111111111111111, 18'b000000000000111101, 18'b111111111111111101, 18'b111111111111101011, 18'b000000000000000000, 18'b000000000000010000, 18'b111111111111100111, 18'b000000000000110010, 18'b000000000000010000, 18'b111111111011010110, 18'b111111111111000101, 18'b000000000000101110, 18'b111111111111111111, 18'b111111111011111101, 18'b111111111110111111, 18'b111111111111110100, 18'b111111111111111111, 18'b111111111111100010, 18'b000000000000000000, 18'b111111111111101011}, 
{18'b000000000000000000, 18'b111111111111111111, 18'b111111111111010001, 18'b111111111110101001, 18'b000000000000010101, 18'b000000000000000000, 18'b000000000000110000, 18'b111111111111111101, 18'b000000000001111111, 18'b111111111111111101, 18'b000000000000000000, 18'b111111111101010000, 18'b111111111111111111, 18'b000000000001000000, 18'b111111111111111111, 18'b111111111101111010, 18'b000000000000000000, 18'b111111111111111010, 18'b000000000010000110, 18'b111111111111111111, 18'b111111111100100000, 18'b111111111111111111, 18'b000000000010000100, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000001000111, 18'b111111111111001111, 18'b000000000000100011, 18'b000000000000000000, 18'b111111111110011000, 18'b000000000000000000, 18'b000000000000000001}, 
{18'b111111111110010001, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111111111100, 18'b000000000011111101, 18'b111111111111000000, 18'b111111111111111101, 18'b111111111111111100, 18'b111111111111101001, 18'b111111111111100110, 18'b000000000000100001, 18'b000000000001000100, 18'b111111111111101101, 18'b000000000001111111, 18'b000000000000000000, 18'b111111111111111111, 18'b111111111101101110, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111111010111, 18'b000000000000000001, 18'b000000000000010011, 18'b000000000000000110, 18'b111111111111111011, 18'b111111111111100101, 18'b111111111110011000, 18'b111111111101101000, 18'b000000000000000000, 18'b111111111111000110, 18'b000000000000010100, 18'b111111111111111111, 18'b000000000000100110}, 
{18'b111111111100101100, 18'b111111111110101111, 18'b111111111110110000, 18'b000000000000000000, 18'b000000000100100100, 18'b111111111110001110, 18'b000000000000000000, 18'b111111111111100100, 18'b111111111100101110, 18'b000000000001000110, 18'b111111111111111111, 18'b000000000100100010, 18'b000000000000000000, 18'b111111111111100111, 18'b111111111111111111, 18'b000000000000010000, 18'b111111111111110110, 18'b000000000000000000, 18'b111111111111101000, 18'b000000000011111101, 18'b000000000000010011, 18'b111111111111101010, 18'b000000000000111000, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111111001110, 18'b111111111111101000, 18'b111111111100010000, 18'b111111111110110110, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111111100001}, 
{18'b000000000001110011, 18'b111111111001100110, 18'b111111111010001101, 18'b111111111110101000, 18'b000000000101010110, 18'b111111111111111111, 18'b111111111101001110, 18'b000000000010000111, 18'b000000000000011110, 18'b000000000000000000, 18'b000000000001101010, 18'b111111111101110101, 18'b000000000000000000, 18'b000000000000000010, 18'b111111111111101111, 18'b000000000000001001, 18'b111111111111001010, 18'b111111111000101000, 18'b000000000001010101, 18'b000000000010110000, 18'b000000000010000111, 18'b000000000000000001, 18'b000000000000001110, 18'b111111111100110001, 18'b111111111010111100, 18'b111111111111111101, 18'b111111111101100110, 18'b111111111100010101, 18'b111111111110011100, 18'b111111111000111110, 18'b000000000011010110, 18'b000000000011011011}, 
{18'b000000000000000000, 18'b000000000000000000, 18'b000000000000000001, 18'b000000000000000000, 18'b000000000010000100, 18'b111111111110100000, 18'b000000000000001001, 18'b000000000000100101, 18'b111111111101001101, 18'b000000000000010010, 18'b111111111111111101, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000001111010, 18'b000000000000011010, 18'b000000000000001011, 18'b000000000000011111, 18'b000000000010101010, 18'b111111111110010000, 18'b000000000000000000, 18'b111111111110101011, 18'b111111111111111111, 18'b000000000010100001, 18'b000000000000000100, 18'b111111111111111110, 18'b111111111011100000, 18'b111111111111111011, 18'b111111111110110000, 18'b111111111111100000, 18'b000000000000000001, 18'b000000000001000101, 18'b000000000000110101}, 
{18'b111111111111101001, 18'b000000000001000100, 18'b111111111101100100, 18'b000000000000001010, 18'b000000000001100011, 18'b111111111111101011, 18'b111111111111111101, 18'b000000000001010011, 18'b000000000000000000, 18'b111111111111111111, 18'b111111111111011110, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111111101110, 18'b111111111111000001, 18'b111111111111011110, 18'b111111111111100011, 18'b111111111111011111, 18'b111111111111000111, 18'b000000000000000000, 18'b111111111111111111, 18'b111111111111101001, 18'b111111111111011101, 18'b000000000011001011, 18'b000000000000000000, 18'b111111111101000111, 18'b111111111111111011, 18'b000000000000111111, 18'b000000000000000000, 18'b000000000000000000, 18'b000000000010000000, 18'b111111111111111111}, 
{18'b111111111111111111, 18'b000000000000000010, 18'b111111111111111111, 18'b111111111110110000, 18'b111111111001000111, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111111111100, 18'b111111111011001101, 18'b000000000000101001, 18'b111111111111001101, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111101000010, 18'b111111111111101000, 18'b111111111111111111, 18'b000000000000000000, 18'b000000000000000100, 18'b000000000000010010, 18'b000000000010110000, 18'b111111111111000010, 18'b111111111101100110, 18'b000000000000000000, 18'b111111111101111011, 18'b111111111111001101, 18'b111111111110001001, 18'b111111111111111100, 18'b111111111111111001, 18'b111111111111110110, 18'b111111111100001110, 18'b111111111111101110, 18'b000000000001111100}, 
{18'b000000000000111001, 18'b000000000001110000, 18'b111111111111111110, 18'b000000000001010001, 18'b111111111110010100, 18'b111111111111000000, 18'b000000000000110000, 18'b000000000000100011, 18'b111111111111100111, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111101011011, 18'b111111111111111111, 18'b000000000001001001, 18'b111111111111000101, 18'b000000000000010001, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000001101010, 18'b111111111101011000, 18'b000000000010001111, 18'b000000000000011000, 18'b000000000000000000, 18'b000000000001101100, 18'b000000000000000001, 18'b111111111111101101, 18'b111111111100111101, 18'b111111111111000111, 18'b111111111110101000, 18'b000000000001011010}, 
{18'b000000000000000000, 18'b000000000000000011, 18'b111111111101000100, 18'b111111111111111110, 18'b000000000001101001, 18'b111111111110110111, 18'b111111111111111001, 18'b111111111111111111, 18'b000000000000001010, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111110010111, 18'b000000000000110001, 18'b000000000000000011, 18'b000000000000000000, 18'b000000000000010011, 18'b111111111111111111, 18'b111111111110110011, 18'b000000000000001001, 18'b000000000000000000, 18'b111111111111101110, 18'b111111111111110100, 18'b000000000010010111, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111101101010, 18'b111111111101011000, 18'b000000000001111011, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000000001110, 18'b000000000010010000}, 
{18'b111111111101010001, 18'b111111111111111111, 18'b111111111110010011, 18'b000000000000000010, 18'b111111111101001011, 18'b000000000000000000, 18'b111111111111111111, 18'b111111111111011110, 18'b111111111011101111, 18'b111111111111110010, 18'b000000000000000000, 18'b111111111111111011, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111111111011, 18'b111111111111100110, 18'b111111111110110100, 18'b111111111111001111, 18'b000000000000100001, 18'b111111111111111110, 18'b111111111111110011, 18'b000000000000000000, 18'b000000000010101100, 18'b111111111111111111, 18'b000000000001001100, 18'b000000000000101110, 18'b111111111110111001, 18'b000000000001101101, 18'b111111111111101000, 18'b000000000000000000, 18'b111111111111111111, 18'b000000000100101010}, 
{18'b111111111101011111, 18'b000000000000001111, 18'b000000000000011001, 18'b111111111111110001, 18'b000000000001111101, 18'b111111111101100101, 18'b111111111111111100, 18'b000000000010000111, 18'b000000000001010001, 18'b000000000000000100, 18'b111111111111111111, 18'b111111111111011100, 18'b111111111111010010, 18'b111111111111011110, 18'b111111111111100110, 18'b000000000000101110, 18'b111111111111111111, 18'b000000000000000100, 18'b000000000001001000, 18'b000000000000000000, 18'b000000000000000000, 18'b000000000000000111, 18'b000000000010000001, 18'b000000000000010111, 18'b000000000000000011, 18'b111111111111001000, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111111111000, 18'b111111111111111001, 18'b111111111111111111, 18'b000000000000100010}, 
{18'b111111111111111111, 18'b000000000000000001, 18'b111111111110010011, 18'b111111111111011001, 18'b000000000010010000, 18'b111111111111111111, 18'b111111111111011000, 18'b000000000001111101, 18'b111111111111100100, 18'b000000000010010101, 18'b000000000000101011, 18'b111111111111000010, 18'b000000000000000000, 18'b000000000000000001, 18'b111111111111111000, 18'b000000000000001010, 18'b111111111111011000, 18'b111111111101111001, 18'b000000000010001110, 18'b000000000001001111, 18'b000000000101000100, 18'b000000000001100110, 18'b000000000001111111, 18'b111111111111111111, 18'b000000000000000000, 18'b000000000000000000, 18'b000000000000011101, 18'b000000000000101000, 18'b111111111100101000, 18'b111111111111111111, 18'b111111111111111101, 18'b111111111111111100}, 
{18'b000000000000000000, 18'b111111111111010011, 18'b111111111111001010, 18'b000000000000000000, 18'b111111111110000011, 18'b000000000000000000, 18'b000000000001100010, 18'b000000000000110111, 18'b000000000000011011, 18'b111111111111001101, 18'b000000000000000000, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111111101010, 18'b000000000001100111, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111101100101, 18'b000000000000000000, 18'b111111111110011101, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111111111101, 18'b000000000000000111, 18'b000000000000001000, 18'b000000000000001110, 18'b000000000001000110, 18'b111111111111011110, 18'b111111111111111100, 18'b111111111100011010, 18'b000000000000101000}, 
{18'b000000000011100010, 18'b111111111111111011, 18'b000000000000100001, 18'b111111111111001010, 18'b111111111111010100, 18'b000000000000010001, 18'b000000000001010010, 18'b000000000000000000, 18'b000000000100001101, 18'b000000000000000000, 18'b111111111111110101, 18'b000000000000001001, 18'b000000000000110000, 18'b111111111111111110, 18'b000000000000011011, 18'b000000000000110100, 18'b111111111111111101, 18'b111111111100011100, 18'b111111111111100011, 18'b111111111111111111, 18'b000000000000111011, 18'b000000000000000000, 18'b111111111111111111, 18'b000000000000111001, 18'b000000000000001001, 18'b111111111101111001, 18'b111111111111001011, 18'b000000000001000011, 18'b111111111111110001, 18'b000000000010000100, 18'b111111111111111111, 18'b111111111110100100}, 
{18'b000000000000000110, 18'b000000000000110100, 18'b111111111111111111, 18'b111111111111101100, 18'b111111111101001011, 18'b111111111111111111, 18'b000000000000010111, 18'b111111111111101000, 18'b000000000001010100, 18'b111111111111101110, 18'b111111111111111111, 18'b111111111111101110, 18'b111111111111111111, 18'b111111111111101101, 18'b000000000000000000, 18'b000000000010100000, 18'b000000000000000000, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000000010001, 18'b000000000001000000, 18'b000000000000000000, 18'b000000000000000010, 18'b000000000000010000, 18'b111111111111111111, 18'b000000000000000000, 18'b000000000000001010, 18'b000000000000000000, 18'b000000000000110001}, 
{18'b111111111101100001, 18'b000000000001000010, 18'b000000000000001001, 18'b111111111111001010, 18'b111111111100110011, 18'b111111111111110110, 18'b000000000000100010, 18'b111111111100110100, 18'b000000000100000101, 18'b000000000000100100, 18'b000000000000001000, 18'b000000000000110000, 18'b000000000000010110, 18'b000000000000000000, 18'b000000000011010000, 18'b111111111111010100, 18'b000000000000000010, 18'b000000000000000000, 18'b111111111111111100, 18'b000000000000000001, 18'b111111111100100010, 18'b000000000000001000, 18'b000000000001001110, 18'b000000000000010011, 18'b000000000000010010, 18'b111111111010101111, 18'b111111111101010001, 18'b111111111110000100, 18'b000000000000000001, 18'b111111111111111111, 18'b000000000010100110, 18'b111111111110010111}, 
{18'b111111111111111001, 18'b111111111110011100, 18'b111111111111001011, 18'b111111111100101110, 18'b111111111101111010, 18'b000000000010101100, 18'b000000000010011110, 18'b111111111110101000, 18'b000000000000010101, 18'b111111111111101100, 18'b111111111111001111, 18'b111111111101111111, 18'b000000000000110100, 18'b111111111101101110, 18'b000000000001100000, 18'b111111111111111111, 18'b000000000010101011, 18'b111111111111111111, 18'b111111111111111100, 18'b111111111110111010, 18'b111111111111101010, 18'b111111111111011110, 18'b111111111101110111, 18'b000000000000101010, 18'b111111111111111111, 18'b111111111111111100, 18'b111111111110001011, 18'b000000000010100001, 18'b000000000010001110, 18'b111111111111010001, 18'b111111111010111101, 18'b000000000001001001}, 
{18'b000000000000000000, 18'b111111111111110010, 18'b111111111111111111, 18'b111111111111001110, 18'b000000000000001110, 18'b000000000000000100, 18'b000000000000100011, 18'b000000000000000010, 18'b000000000000111100, 18'b111111111111111111, 18'b000000000000000000, 18'b000000000000110000, 18'b000000000000000000, 18'b000000000000000110, 18'b111111111110111100, 18'b111111111111001000, 18'b000000000000000000, 18'b000000000001011101, 18'b000000000000011101, 18'b000000000001000000, 18'b111111111111110111, 18'b111111111110101110, 18'b111111111111111111, 18'b000000000000100110, 18'b111111111111111111, 18'b000000000000010000, 18'b111111111111111101, 18'b000000000000100010, 18'b000000000000000000, 18'b000000000000101010, 18'b111111111100111101, 18'b111111111111111111}, 
{18'b000000000010011110, 18'b111111111111111011, 18'b000000000001001100, 18'b111111111101100011, 18'b111111111110011101, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000000001110, 18'b000000000000000001, 18'b111111111110111111, 18'b000000000000000000, 18'b000000000000000001, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111110111101, 18'b000000000001001001, 18'b111111111111111111, 18'b111111111111110000, 18'b000000000000000000, 18'b000000000000111101, 18'b111111111110011001, 18'b000000000000111011, 18'b000000000001000111, 18'b000000000001000010, 18'b111111111111111111, 18'b000000000100011010, 18'b111111111110110001, 18'b000000000010111010, 18'b111111111111100101, 18'b111111111101000111, 18'b111111111110100111, 18'b000000000001000111}, 
{18'b111111111011101001, 18'b111111111111110010, 18'b111111111110110001, 18'b111111111111111111, 18'b000000000010000101, 18'b111111111110100100, 18'b111111111111100001, 18'b000000000001111001, 18'b000000000000110000, 18'b111111111110000110, 18'b000000000000000000, 18'b111111111111110001, 18'b111111111111111010, 18'b000000000001000110, 18'b111111111110000010, 18'b111111111111111010, 18'b000000000000000000, 18'b111111111111111111, 18'b111111111111110111, 18'b000000000000000000, 18'b111111111110011110, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111101010111, 18'b000000000000100011, 18'b000000000100111101, 18'b000000000010110001, 18'b111111111111101101, 18'b111111111110101101, 18'b111111111100011010, 18'b000000000000000000, 18'b111111111111100111}, 
{18'b000000000000001010, 18'b000000000001101101, 18'b000000000000001010, 18'b111111111110110010, 18'b000000000000000010, 18'b111111111111110010, 18'b000000000000000000, 18'b000000000001101010, 18'b000000000001101110, 18'b111111111110111011, 18'b000000000001000111, 18'b000000000000001100, 18'b111111111111111111, 18'b111111111111111000, 18'b111111111110101110, 18'b000000000010000001, 18'b111111111111101010, 18'b111111111101011010, 18'b000000000000111010, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000000111011, 18'b111111111111011001, 18'b111111111111111101, 18'b111111111111100101, 18'b000000000000101101, 18'b111111111110111000, 18'b000000000001000100, 18'b111111111101000101, 18'b000000000000101001, 18'b111111111111111111, 18'b000000000001010000}, 
{18'b111111111111101010, 18'b000000000000000000, 18'b000000000000101101, 18'b000000000000000000, 18'b111111111111100000, 18'b111111111111111110, 18'b000000000000110100, 18'b111111111111111111, 18'b000000000000000000, 18'b000000000000000010, 18'b000000000000000000, 18'b000000000000001010, 18'b111111111111001001, 18'b000000000000000101, 18'b000000000000111000, 18'b000000000000010111, 18'b000000000000110110, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000001000001, 18'b000000000001111110, 18'b111111111111001101, 18'b000000000000000000, 18'b111111111111111110, 18'b000000000000000101, 18'b111111111100010011, 18'b111111111111111111, 18'b111111111111011011, 18'b111111111111111111, 18'b000000000100100001, 18'b000000000000000000, 18'b111111111110010110}, 
{18'b111111111111110010, 18'b111111111111000010, 18'b111111111111111011, 18'b000000000000000011, 18'b000000000000101110, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111111110100, 18'b000000000000100100, 18'b111111111111111011, 18'b000000000000000000, 18'b000000000000010000, 18'b000000000010010111, 18'b111111111111001011, 18'b000000000000000110, 18'b111111111001001101, 18'b111111111111111010, 18'b111111111111100001, 18'b000000000000000100, 18'b111111111111100110, 18'b000000000000101111, 18'b111111111110001101, 18'b000000000000111010, 18'b000000000000110101, 18'b111111111111111001, 18'b111111111010010011, 18'b111111111110001010, 18'b111111111111110100, 18'b111111111111110110, 18'b000000000011000111, 18'b111111111111111101, 18'b000000000001001110}, 
{18'b000000000000011000, 18'b000000000000000000, 18'b000000000001011001, 18'b111111111111000101, 18'b111111111111011100, 18'b000000000001111001, 18'b111111111110101110, 18'b000000000000011101, 18'b111111111101100001, 18'b000000000000000100, 18'b000000000000001000, 18'b111111111111010101, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111110011111, 18'b000000000011011101, 18'b111111111110000001, 18'b111111111111111001, 18'b000000000000111100, 18'b111111111111111111, 18'b000000000000100011, 18'b111111111100001010, 18'b000000000010100000, 18'b111111111111111111, 18'b111111111111000000, 18'b000000000011111000, 18'b000000000001001010, 18'b111111111110101111, 18'b111111111110111011, 18'b111111111011101100, 18'b111111111111111010, 18'b000000000000001000}, 
{18'b111111111111111111, 18'b000000000000000011, 18'b111111111111101110, 18'b111111111101110110, 18'b111111111111111111, 18'b111111111100110111, 18'b000000000000000000, 18'b000000000010011011, 18'b000000000001111101, 18'b000000000000001001, 18'b000000000000000000, 18'b111111111111000111, 18'b000000000010101010, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000011011110, 18'b000000000000000000, 18'b111111111111101011, 18'b111111111111100101, 18'b111111111101011011, 18'b000000000001000011, 18'b000000000000000000, 18'b000000000000000000, 18'b000000000000010000, 18'b111111111111011011, 18'b111111111100010100, 18'b000000000010001101, 18'b111111111100011100, 18'b000000000000011010, 18'b111111111111010111, 18'b000000000000000000}, 
{18'b000000000000011111, 18'b000000000001011111, 18'b000000000000000100, 18'b111111111111111110, 18'b111111111100010100, 18'b000000000000000000, 18'b111111111111111111, 18'b000000000001111100, 18'b000000000010001101, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000000000000, 18'b000000000000000001, 18'b000000000000000000, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111111111111, 18'b000000000001010111, 18'b111111111111001011, 18'b111111111100100010, 18'b111111111111101111, 18'b111111111111001101, 18'b111111111111001111, 18'b111111111111011100, 18'b111111111111111111, 18'b111111111111011111, 18'b111111111111110100, 18'b111111111111111010, 18'b000000000001001000, 18'b111111111111111111, 18'b000000000011101101}
};

localparam logic signed [17:0] bias [32] = '{
18'b000000001011110010,  // 1.474280834197998
18'b000000000101100010,  // 0.6914801001548767
18'b000000001011100001,  // 1.4406442642211914
18'b000000001011010000,  // 1.408045768737793
18'b000000000111111001,  // 0.9864811301231384
18'b000000000110111010,  // 0.8636202812194824
18'b111111111011000100,  // -0.6153604388237
18'b000000000011110111,  // 0.4839226007461548
18'b000000000011111000,  // 0.4862793982028961
18'b000000000010111110,  // 0.37162142992019653
18'b000000000011101011,  // 0.45989668369293213
18'b000000001010011001,  // 1.2998151779174805
18'b111111110111110111,  // -1.016528844833374
18'b111111111101001011,  // -0.35249894857406616
18'b000000000011100100,  // 0.44582197070121765
18'b111111111111000110,  // -0.1119980737566948
18'b111111111111011101,  // -0.06717441976070404
18'b000000000000000010,  // 0.00487547367811203
18'b000000000001100011,  // 0.1946917623281479
18'b111111111001110000,  // -0.7796769738197327
18'b000000000101110101,  // 0.7287401556968689
18'b000000001101101110,  // 1.714877724647522
18'b111111110011001110,  // -1.5971007347106934
18'b000000000000100101,  // 0.07393483817577362
18'b000000000010100101,  // 0.3225609362125397
18'b000000000110110000,  // 0.8453295230865479
18'b000000000111001100,  // 0.898597240447998
18'b000000000010000010,  // 0.2548799514770508
18'b000000000111110010,  // 0.9735668301582336
18'b000000001001000000,  // 1.1261906623840332
18'b000000000011100101,  // 0.44768181443214417
18'b111111101101000011   // -2.3676068782806396
};
endpackage