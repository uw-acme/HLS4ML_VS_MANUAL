//Width: 4
//Int: 2
package dense_3_gen;

localparam logic signed [3:0] weights [32][32] = '{
{4'b1111, 4'b1110, 4'b1110, 4'b1111, 4'b0001, 4'b0000, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b1110, 4'b1111, 4'b0011, 4'b1111, 4'b1100, 4'b1111, 4'b0000, 4'b0010, 4'b1111, 4'b1100, 4'b1111, 4'b0000, 4'b1110, 4'b0000, 4'b0100, 4'b1010, 4'b1111, 4'b1110, 4'b1111, 4'b0010, 4'b1111},
{4'b0011, 4'b0111, 4'b0010, 4'b1101, 4'b0001, 4'b1111, 4'b1111, 4'b0100, 4'b0000, 4'b1111, 4'b1111, 4'b1110, 4'b1111, 4'b0010, 4'b1000, 4'b1110, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b0000, 4'b1111, 4'b1111, 4'b1100, 4'b0000, 4'b0010, 4'b1111, 4'b1101, 4'b0000, 4'b0000},
{4'b1100, 4'b0001, 4'b0000, 4'b0001, 4'b1101, 4'b0000, 4'b0000, 4'b1101, 4'b0010, 4'b1111, 4'b1111, 4'b1010, 4'b1111, 4'b0010, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b1101, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0100, 4'b0000, 4'b1101, 4'b0011, 4'b0000, 4'b0001, 4'b1111, 4'b0000, 4'b0111},
{4'b0011, 4'b1111, 4'b1111, 4'b0101, 4'b0101, 4'b0000, 4'b0000, 4'b0011, 4'b1110, 4'b1111, 4'b1101, 4'b0000, 4'b0001, 4'b1101, 4'b0000, 4'b1111, 4'b1111, 4'b1111, 4'b0000, 4'b0000, 4'b0000, 4'b1111, 4'b0101, 4'b0011, 4'b0011, 4'b0010, 4'b0011, 4'b0000, 4'b1111, 4'b0100, 4'b0010, 4'b1111},
{4'b0100, 4'b1111, 4'b1101, 4'b1010, 4'b0100, 4'b0000, 4'b1101, 4'b1110, 4'b1111, 4'b1010, 4'b1111, 4'b0100, 4'b0101, 4'b0100, 4'b1011, 4'b1010, 4'b0000, 4'b1111, 4'b0010, 4'b0001, 4'b1110, 4'b1111, 4'b0110, 4'b0111, 4'b0001, 4'b1011, 4'b0001, 4'b1110, 4'b1110, 4'b1111, 4'b0001, 4'b0101},
{4'b0000, 4'b1111, 4'b1110, 4'b1110, 4'b0011, 4'b0000, 4'b1110, 4'b1111, 4'b1101, 4'b1111, 4'b1111, 4'b0001, 4'b0000, 4'b0011, 4'b1100, 4'b1111, 4'b0001, 4'b1110, 4'b1110, 4'b1111, 4'b0000, 4'b0010, 4'b0100, 4'b1111, 4'b1111, 4'b0011, 4'b1100, 4'b1111, 4'b1110, 4'b1111, 4'b1111, 4'b0000},
{4'b0001, 4'b1101, 4'b0001, 4'b1111, 4'b1111, 4'b0001, 4'b1111, 4'b1011, 4'b1111, 4'b1110, 4'b1100, 4'b0100, 4'b0000, 4'b0101, 4'b0111, 4'b0000, 4'b1111, 4'b1101, 4'b1111, 4'b0010, 4'b1010, 4'b0001, 4'b0011, 4'b0000, 4'b0001, 4'b0111, 4'b1101, 4'b1111, 4'b1110, 4'b0100, 4'b1111, 4'b1111},
{4'b1011, 4'b0000, 4'b1011, 4'b0011, 4'b0000, 4'b0001, 4'b0000, 4'b0000, 4'b1111, 4'b0001, 4'b0111, 4'b1111, 4'b0011, 4'b0101, 4'b0110, 4'b0000, 4'b0000, 4'b1100, 4'b0011, 4'b1111, 4'b1011, 4'b1110, 4'b0000, 4'b1111, 4'b1100, 4'b0111, 4'b1110, 4'b0000, 4'b0000, 4'b0111, 4'b0001, 4'b0011},
{4'b0011, 4'b1111, 4'b0000, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b0001, 4'b0010, 4'b1110, 4'b0001, 4'b0001, 4'b0000, 4'b0011, 4'b1110, 4'b1010, 4'b0000, 4'b1111, 4'b1111, 4'b1100, 4'b1111, 4'b0000, 4'b1110, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1111, 4'b0000, 4'b1101},
{4'b1111, 4'b0011, 4'b0000, 4'b0000, 4'b0110, 4'b0011, 4'b1111, 4'b1100, 4'b0001, 4'b1010, 4'b0111, 4'b1111, 4'b0000, 4'b0011, 4'b0001, 4'b0000, 4'b1101, 4'b0000, 4'b0000, 4'b0000, 4'b0010, 4'b1111, 4'b1101, 4'b0000, 4'b1111, 4'b0111, 4'b0011, 4'b1111, 4'b1111, 4'b0101, 4'b1111, 4'b1111},
{4'b1100, 4'b0001, 4'b1111, 4'b1111, 4'b1110, 4'b1101, 4'b0000, 4'b0001, 4'b1111, 4'b1111, 4'b1011, 4'b0010, 4'b0010, 4'b0000, 4'b0111, 4'b1100, 4'b0001, 4'b1101, 4'b0010, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b0000, 4'b1100, 4'b0000, 4'b1100, 4'b1111, 4'b1111, 4'b0101, 4'b1110, 4'b0000},
{4'b1111, 4'b0001, 4'b0000, 4'b0011, 4'b1111, 4'b1111, 4'b0000, 4'b1111, 4'b1111, 4'b0101, 4'b0110, 4'b0000, 4'b1101, 4'b1010, 4'b1111, 4'b0000, 4'b0000, 4'b1111, 4'b1100, 4'b0011, 4'b0000, 4'b0011, 4'b1111, 4'b0100, 4'b0001, 4'b0010, 4'b0100, 4'b1111, 4'b1101, 4'b1100, 4'b1111, 4'b1011},
{4'b1110, 4'b1111, 4'b0001, 4'b1101, 4'b0001, 4'b1111, 4'b1110, 4'b1111, 4'b1111, 4'b0000, 4'b0001, 4'b1111, 4'b0000, 4'b0010, 4'b1011, 4'b1110, 4'b0010, 4'b1111, 4'b0000, 4'b1111, 4'b0010, 4'b0000, 4'b1111, 4'b0000, 4'b0010, 4'b1111, 4'b0000, 4'b1100, 4'b1110, 4'b1111, 4'b0001, 4'b0000},
{4'b1100, 4'b0011, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b1111, 4'b0110, 4'b1111, 4'b1111, 4'b0010, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0011, 4'b0001, 4'b0001, 4'b1111, 4'b0010, 4'b0001, 4'b0000, 4'b1111, 4'b0010, 4'b1111, 4'b1101, 4'b1111, 4'b1111, 4'b0001, 4'b0000, 4'b0010, 4'b0100},
{4'b1111, 4'b1101, 4'b0000, 4'b1111, 4'b0111, 4'b1110, 4'b1011, 4'b0000, 4'b0000, 4'b1111, 4'b0000, 4'b0011, 4'b0011, 4'b0000, 4'b0000, 4'b1111, 4'b0000, 4'b1111, 4'b0000, 4'b0001, 4'b1111, 4'b0000, 4'b0010, 4'b0000, 4'b1111, 4'b1101, 4'b0010, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111},
{4'b0000, 4'b1111, 4'b1111, 4'b1110, 4'b1100, 4'b0101, 4'b0000, 4'b0001, 4'b0010, 4'b0000, 4'b1111, 4'b0100, 4'b0010, 4'b1101, 4'b1111, 4'b1111, 4'b1101, 4'b1111, 4'b0000, 4'b1111, 4'b0001, 4'b1111, 4'b0000, 4'b0001, 4'b1111, 4'b1101, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b1101, 4'b0000},
{4'b1110, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b0001, 4'b1111, 4'b0000, 4'b0001, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b1111, 4'b0100, 4'b1111, 4'b0010, 4'b1111, 4'b0001, 4'b0001, 4'b0001, 4'b0000, 4'b1111, 4'b1110, 4'b1110, 4'b0001, 4'b1111, 4'b0000, 4'b1111, 4'b0010},
{4'b1111, 4'b1101, 4'b1101, 4'b1111, 4'b0101, 4'b1111, 4'b0000, 4'b0100, 4'b1111, 4'b0000, 4'b1101, 4'b1100, 4'b0100, 4'b0001, 4'b1111, 4'b1110, 4'b0001, 4'b0000, 4'b1110, 4'b0000, 4'b0001, 4'b1111, 4'b0010, 4'b1000, 4'b0000, 4'b0010, 4'b1111, 4'b0000, 4'b1110, 4'b1111, 4'b1110, 4'b1111},
{4'b0010, 4'b0011, 4'b0100, 4'b1110, 4'b0011, 4'b0010, 4'b0000, 4'b0100, 4'b0011, 4'b1111, 4'b0110, 4'b1101, 4'b0101, 4'b0100, 4'b1111, 4'b1111, 4'b0000, 4'b0000, 4'b0010, 4'b1100, 4'b0010, 4'b1110, 4'b1100, 4'b1111, 4'b0011, 4'b1011, 4'b1101, 4'b1111, 4'b1111, 4'b1011, 4'b0011, 4'b0000},
{4'b1111, 4'b0000, 4'b1111, 4'b1111, 4'b1101, 4'b0000, 4'b0000, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b1111, 4'b0001, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b0100, 4'b1101, 4'b0000, 4'b1111, 4'b0001, 4'b0010, 4'b1111, 4'b1110, 4'b0000, 4'b0111, 4'b1111, 4'b1111, 4'b0011, 4'b0000, 4'b0111},
{4'b1100, 4'b0000, 4'b1110, 4'b0011, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b1110, 4'b1111, 4'b0000, 4'b1100, 4'b0000, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b0000, 4'b0000, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b1111, 4'b0000, 4'b0000, 4'b0101, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b1111},
{4'b1111, 4'b1111, 4'b0010, 4'b0000, 4'b1101, 4'b0000, 4'b0010, 4'b1111, 4'b0000, 4'b1111, 4'b0001, 4'b0000, 4'b0011, 4'b1100, 4'b1111, 4'b1111, 4'b0010, 4'b1101, 4'b0000, 4'b1010, 4'b1111, 4'b1111, 4'b1111, 4'b0010, 4'b1111, 4'b1110, 4'b0001, 4'b0000, 4'b0011, 4'b0100, 4'b1101, 4'b1100},
{4'b0001, 4'b0000, 4'b1101, 4'b1111, 4'b1111, 4'b0000, 4'b0001, 4'b0011, 4'b0000, 4'b0000, 4'b0001, 4'b1100, 4'b1111, 4'b1011, 4'b0100, 4'b0000, 4'b1111, 4'b1011, 4'b1111, 4'b1111, 4'b1111, 4'b0000, 4'b0000, 4'b1111, 4'b0000, 4'b0011, 4'b0011, 4'b0011, 4'b0010, 4'b0000, 4'b0001, 4'b0110},
{4'b1111, 4'b1110, 4'b0011, 4'b1111, 4'b0001, 4'b0001, 4'b1111, 4'b1110, 4'b1111, 4'b1011, 4'b0100, 4'b0000, 4'b0011, 4'b0101, 4'b1111, 4'b1001, 4'b1111, 4'b0100, 4'b1110, 4'b1110, 4'b0000, 4'b0000, 4'b1100, 4'b1110, 4'b1111, 4'b1111, 4'b0001, 4'b0110, 4'b0010, 4'b1111, 4'b0001, 4'b0000},
{4'b0000, 4'b0100, 4'b0000, 4'b0010, 4'b0111, 4'b1111, 4'b1111, 4'b1111, 4'b0010, 4'b1110, 4'b1111, 4'b0011, 4'b0000, 4'b0000, 4'b0111, 4'b1111, 4'b0000, 4'b0010, 4'b1111, 4'b0010, 4'b1111, 4'b1111, 4'b1100, 4'b0001, 4'b0010, 4'b1111, 4'b1111, 4'b0000, 4'b0100, 4'b1010, 4'b0000, 4'b1111},
{4'b0000, 4'b1101, 4'b0000, 4'b1111, 4'b0000, 4'b0100, 4'b1010, 4'b0000, 4'b0011, 4'b1101, 4'b1111, 4'b0000, 4'b1111, 4'b0001, 4'b0001, 4'b1111, 4'b0001, 4'b0000, 4'b0000, 4'b0011, 4'b1111, 4'b1100, 4'b1011, 4'b1110, 4'b1011, 4'b0010, 4'b0101, 4'b0011, 4'b1111, 4'b1101, 4'b1110, 4'b0000},
{4'b0000, 4'b1100, 4'b1111, 4'b0001, 4'b1100, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0000, 4'b0010, 4'b1111, 4'b0000, 4'b0000, 4'b0001, 4'b1111, 4'b0000, 4'b1111, 4'b1101, 4'b1100, 4'b1111, 4'b1100, 4'b1110, 4'b1101, 4'b0111, 4'b0000, 4'b1111, 4'b0011, 4'b0111, 4'b0011, 4'b1000, 4'b1111},
{4'b0011, 4'b1111, 4'b0010, 4'b1111, 4'b0100, 4'b1111, 4'b0001, 4'b0011, 4'b0010, 4'b1100, 4'b1111, 4'b0001, 4'b0001, 4'b1111, 4'b0001, 4'b0000, 4'b0011, 4'b0000, 4'b0011, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b0010, 4'b1110, 4'b1111, 4'b0000, 4'b0000, 4'b0000, 4'b0010, 4'b1101, 4'b1111},
{4'b1111, 4'b1111, 4'b1100, 4'b0010, 4'b0010, 4'b1111, 4'b1111, 4'b1110, 4'b0000, 4'b1111, 4'b1110, 4'b1110, 4'b0100, 4'b0000, 4'b1111, 4'b1111, 4'b0010, 4'b1111, 4'b1111, 4'b1110, 4'b0011, 4'b0000, 4'b0001, 4'b1111, 4'b0001, 4'b0000, 4'b0000, 4'b0010, 4'b1110, 4'b1111, 4'b0001, 4'b1111},
{4'b1111, 4'b1110, 4'b0101, 4'b1111, 4'b0010, 4'b1110, 4'b0000, 4'b0000, 4'b1100, 4'b1111, 4'b1111, 4'b0000, 4'b1101, 4'b0001, 4'b0010, 4'b0001, 4'b0001, 4'b1111, 4'b1010, 4'b1111, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b0010, 4'b1111, 4'b1111, 4'b0011, 4'b1101, 4'b1110, 4'b0011, 4'b0000},
{4'b0011, 4'b0010, 4'b0000, 4'b1111, 4'b1111, 4'b1111, 4'b0000, 4'b1111, 4'b1111, 4'b1111, 4'b0000, 4'b0001, 4'b0000, 4'b0000, 4'b1111, 4'b0000, 4'b1111, 4'b0000, 4'b1111, 4'b1111, 4'b0000, 4'b0000, 4'b0001, 4'b0000, 4'b0000, 4'b1011, 4'b1110, 4'b0000, 4'b0000, 4'b0000, 4'b1111, 4'b0000},
{4'b0010, 4'b1000, 4'b1111, 4'b1111, 4'b1110, 4'b1111, 4'b0000, 4'b0100, 4'b1111, 4'b1111, 4'b0001, 4'b1011, 4'b0000, 4'b1100, 4'b0110, 4'b1111, 4'b1110, 4'b1100, 4'b1111, 4'b1010, 4'b1010, 4'b1111, 4'b0000, 4'b0000, 4'b0010, 4'b1111, 4'b1110, 4'b1111, 4'b1111, 4'b0000, 4'b1111, 4'b1010}
};
localparam logic signed [3:0] bias [32] = '{
4'b0010,
4'b0011,
4'b0010,
4'b0010,
4'b0111,
4'b1100,
4'b0111,
4'b1011,
4'b1110,
4'b0111,
4'b0001,
4'b0100,
4'b0111,
4'b1000,
4'b0111,
4'b0111,
4'b1110,
4'b0111,
4'b0011,
4'b0100,
4'b0110,
4'b0011,
4'b0010,
4'b0100,
4'b1111,
4'b1110,
4'b1110,
4'b1011,
4'b0000,
4'b1101,
4'b0100,
4'b1100
};
endpackage