// Width: 17
// NFRAC: 8
package dense_1_17_8;

localparam logic signed [16:0] weights [16][64] = '{ 
{17'b00000000001000001, 17'b11111111101011001, 17'b11111111111010001, 17'b11111111111000110, 17'b11111111110011000, 17'b00000000000011100, 17'b11111111011110110, 17'b00000000000000000, 17'b00000000000001110, 17'b00000000001000011, 17'b00000000000000000, 17'b11111111110011000, 17'b11111111111111111, 17'b00000000000110101, 17'b00000000000001000, 17'b11111111110111101, 17'b00000000000111011, 17'b00000000000001111, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000001100000, 17'b11111111110101011, 17'b11111111111111010, 17'b00000000001111001, 17'b11111111110101101, 17'b11111111101010001, 17'b11111111110111001, 17'b11111111111001110, 17'b11111111111100101, 17'b11111111111111111, 17'b00000000000001001, 17'b00000000000111110, 17'b00000000000110010, 17'b11111111111111100, 17'b00000000000000000, 17'b00000000001001111, 17'b11111111111111011, 17'b11111111110111111, 17'b00000000000000110, 17'b00000000000110001, 17'b11111111111111100, 17'b00000000001000110, 17'b11111111110111011, 17'b00000000011101101, 17'b11111111111111111, 17'b00000000001110011, 17'b00000000000000000, 17'b00000000000101111, 17'b00000000000110010, 17'b11111111111111001, 17'b00000000000000000, 17'b00000000000101001, 17'b00000000000110111, 17'b00000000000010011, 17'b11111111111100010, 17'b11111111110110000, 17'b00000000010001001, 17'b11111111110000000, 17'b00000000001110111, 17'b11111111110100101, 17'b00000000011001011, 17'b11111111111111110, 17'b00000000000000010, 17'b00000000000010100}, 
{17'b00000000000000000, 17'b11111111110101101, 17'b11111111111011110, 17'b11111111110111000, 17'b11111111110101110, 17'b00000000000011011, 17'b11111111100111110, 17'b11111111111111111, 17'b11111111111000101, 17'b00000000000101100, 17'b00000000000000001, 17'b11111111111101001, 17'b00000000000110010, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000000110101, 17'b11111111111111110, 17'b00000000000000000, 17'b11111111111010001, 17'b11111111110111111, 17'b00000000001110001, 17'b11111111111101011, 17'b00000000000001100, 17'b00000000010110010, 17'b00000000001000001, 17'b11111111111000101, 17'b11111111111000100, 17'b11111111111111111, 17'b11111111111100110, 17'b11111111110011000, 17'b11111111111110000, 17'b00000000001110100, 17'b00000000001000111, 17'b00000000010001100, 17'b00000000010100001, 17'b00000000000001100, 17'b11111111111100001, 17'b11111111110010000, 17'b00000000000001110, 17'b00000000000110000, 17'b00000000000000101, 17'b00000000000110100, 17'b11111111111001001, 17'b00000000001000000, 17'b00000000000101100, 17'b00000000000001100, 17'b11111111110101000, 17'b00000000000010100, 17'b00000000001000010, 17'b00000000000000111, 17'b00000000000000110, 17'b00000000100101000, 17'b11111111111101100, 17'b11111111111100110, 17'b11111111111110010, 17'b11111111111111110, 17'b00000000001000001, 17'b11111111110100001, 17'b00000000011111100, 17'b00000000000000001, 17'b00000000010000101, 17'b00000000000111101, 17'b00000000011010010, 17'b00000000000100100}, 
{17'b11111111111111110, 17'b00000000000000000, 17'b11111111111101010, 17'b11111111111010010, 17'b11111111111010000, 17'b00000000000001010, 17'b00000000101111011, 17'b11111111111111111, 17'b11111111010111011, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111111011, 17'b11111111111000101, 17'b00000000000000000, 17'b11111111111111101, 17'b00000000000101011, 17'b00000000011100111, 17'b11111111111111111, 17'b00000000000010010, 17'b00000000000000000, 17'b00000000001101001, 17'b11111111101000111, 17'b00000000010010011, 17'b11111111101001001, 17'b00000000011110010, 17'b11111111110100111, 17'b11111111111000001, 17'b11111111101001000, 17'b00000000101000110, 17'b00000000001000110, 17'b00000000000000010, 17'b00000000010000100, 17'b00000000100000101, 17'b11111111011001110, 17'b11111111111100111, 17'b00000000000001000, 17'b11111111111000100, 17'b00000000011100101, 17'b11111111111110101, 17'b00000000001010000, 17'b00000000001010101, 17'b00000000001011110, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111111011, 17'b00000000000101000, 17'b11111111110111000, 17'b11111111111010100, 17'b11111111111111011, 17'b00000000001100100, 17'b11111111111010010, 17'b00000000000100110, 17'b11111111111111111, 17'b00000000000100010, 17'b11111111111010011, 17'b11111111111111111, 17'b11111111110110001, 17'b11111111101010100, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000110001010, 17'b00000000000000011, 17'b11111111111111111, 17'b11111111110110000}, 
{17'b11111111110001010, 17'b11111111110100001, 17'b11111111101001110, 17'b00000000001001110, 17'b11111111110101111, 17'b11111111010100111, 17'b11111111111100010, 17'b11111111110110001, 17'b00000000000111001, 17'b11111111111111111, 17'b00000000101000011, 17'b11111111111100100, 17'b11111111100110111, 17'b00000000010010100, 17'b00000000000000110, 17'b11111111111111111, 17'b11111111110001110, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111000110, 17'b11111111011011001, 17'b11111111111100011, 17'b11111111101001101, 17'b00000000000110010, 17'b11111111110011100, 17'b11111111100010100, 17'b00000000001010000, 17'b00000000010111100, 17'b00000000101001011, 17'b11111111110001010, 17'b11111111101101010, 17'b00000000000010010, 17'b00000000010000000, 17'b11111111100101000, 17'b11111111110101111, 17'b00000000000000000, 17'b11111111101000110, 17'b00000000000111110, 17'b11111111110001111, 17'b00000000000011110, 17'b00000000001110101, 17'b00000000000101000, 17'b00000000000000000, 17'b00000000000000101, 17'b00000000010001101, 17'b11111111111001100, 17'b11111111111111111, 17'b11111111110100111, 17'b11111111111111111, 17'b11111111111100111, 17'b11111111101100010, 17'b00000000000010110, 17'b11111111111111111, 17'b00000000000110111, 17'b00000000001010000, 17'b00000000010100101, 17'b11111111100001000, 17'b11111111100010010, 17'b11111111101001011, 17'b00000000011011101, 17'b00000000110111111, 17'b11111111100011001, 17'b11111111111110010, 17'b00000000001101111}, 
{17'b00000000001010111, 17'b11111111101100001, 17'b11111111110111101, 17'b11111111111111111, 17'b11111111111011000, 17'b00000000001010111, 17'b00000000000110000, 17'b11111111111111111, 17'b11111111101100111, 17'b11111111111000010, 17'b11111111110100001, 17'b00000000000001101, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111110101, 17'b00000000001011011, 17'b00000000000100010, 17'b11111111110011011, 17'b00000000000000111, 17'b00000000000000011, 17'b00000000000110101, 17'b11111111111100001, 17'b00000000000010011, 17'b11111111111111011, 17'b00000000100010000, 17'b11111111111010000, 17'b11111111110111000, 17'b11111111110011000, 17'b00000000000000000, 17'b00000000000101010, 17'b00000000000011101, 17'b00000000001000110, 17'b11111111111111100, 17'b00000000000010010, 17'b00000000000100001, 17'b11111111111111111, 17'b00000000000000001, 17'b00000000011100001, 17'b11111111110110110, 17'b11111111111101100, 17'b00000000001101110, 17'b00000000000111111, 17'b11111111110000010, 17'b00000000000000001, 17'b11111111011101110, 17'b11111111111111111, 17'b11111111111100000, 17'b00000000000000011, 17'b11111111111111111, 17'b11111111111111001, 17'b11111111111111111, 17'b00000000000110000, 17'b11111111111111110, 17'b00000000001010001, 17'b11111111111001111, 17'b11111111101000011, 17'b11111111110001000, 17'b11111111101111101, 17'b11111111101100010, 17'b00000000010111111, 17'b00000000101011111, 17'b00000000011001010, 17'b00000000000011111, 17'b11111111111111111}, 
{17'b11111111110001101, 17'b11111111101011110, 17'b00000000000000000, 17'b00000000001001110, 17'b00000000001001001, 17'b11111111111001001, 17'b00000000010010101, 17'b11111111111111111, 17'b00000000000111110, 17'b11111111111111111, 17'b11111111111111101, 17'b11111111111101101, 17'b11111111111010010, 17'b00000000010010100, 17'b11111111111101001, 17'b00000000000000000, 17'b11111111101100000, 17'b11111111110100101, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111111110011, 17'b11111111110101111, 17'b11111111110101110, 17'b00000000001110111, 17'b11111111110101110, 17'b11111111111111111, 17'b00000000001000001, 17'b11111111111101101, 17'b11111111100010001, 17'b11111111111111111, 17'b11111111111101110, 17'b11111111111111101, 17'b11111111111111101, 17'b00000000000001010, 17'b00000000000100001, 17'b00000000001011000, 17'b00000000000000011, 17'b11111111111100110, 17'b11111111110111100, 17'b11111111111111111, 17'b11111111111010100, 17'b11111111101111001, 17'b00000000001100110, 17'b00000000000000010, 17'b00000000010011010, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000000011000, 17'b11111111110010100, 17'b00000000000111011, 17'b00000000000000000, 17'b11111111111100110, 17'b11111111110100011, 17'b00000000001100010, 17'b11111111111111111, 17'b00000000001011000, 17'b00000000000110111, 17'b00000000000110100, 17'b11111111111111011, 17'b11111111111111101, 17'b11111111100110001, 17'b11111111111011111, 17'b11111111111110001, 17'b11111111111111111}, 
{17'b11111111110110111, 17'b11111111110101010, 17'b11111111110010001, 17'b11111111111101110, 17'b11111111111011101, 17'b00000000000011010, 17'b11111111101001101, 17'b11111111111011001, 17'b11111111111000110, 17'b11111111111111111, 17'b11111111110110110, 17'b00000000001011001, 17'b00000000000001001, 17'b00000000000100011, 17'b00000000001001111, 17'b00000000000000000, 17'b00000000011001100, 17'b00000000000010110, 17'b00000000000111110, 17'b00000000001000100, 17'b11111111111010111, 17'b00000000001011101, 17'b11111111111000001, 17'b11111111101111111, 17'b00000000000101100, 17'b00000000010000100, 17'b11111111111111110, 17'b00000000000001101, 17'b11111111100001100, 17'b00000000001001001, 17'b00000000001000100, 17'b11111111110100000, 17'b00000000001111000, 17'b00000000010101010, 17'b00000000000000000, 17'b00000000001010111, 17'b11111111111111111, 17'b00000000001001000, 17'b00000000000110010, 17'b00000000000000000, 17'b11111111111100001, 17'b11111111110100010, 17'b00000000000100100, 17'b00000000001111011, 17'b00000000010000100, 17'b11111111111010100, 17'b11111111111101010, 17'b11111111111001111, 17'b11111111111011101, 17'b00000000000011110, 17'b00000000000000000, 17'b00000000000001000, 17'b00000000000000000, 17'b00000000000101110, 17'b11111111111010011, 17'b00000000011000101, 17'b00000000001011011, 17'b11111111111111001, 17'b00000000001100011, 17'b00000000000110111, 17'b11111111001011111, 17'b11111111101101100, 17'b11111111111010011, 17'b11111111111111101}, 
{17'b00000000000000001, 17'b00000000000111101, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111110101101, 17'b11111111111111000, 17'b11111111110111110, 17'b00000000000000000, 17'b00000000000000111, 17'b00000000001100011, 17'b00000000000000011, 17'b11111111110011111, 17'b11111111111101111, 17'b00000000000000000, 17'b11111111111110010, 17'b11111111110001100, 17'b11111111100100110, 17'b11111111111111111, 17'b11111111101100101, 17'b11111111110001101, 17'b11111111110011100, 17'b00000000001011000, 17'b00000000000001100, 17'b11111111111011011, 17'b11111111110010000, 17'b00000000000100111, 17'b00000000000000000, 17'b00000000001111111, 17'b00000000011001110, 17'b11111111111110101, 17'b00000000000000000, 17'b00000000000111011, 17'b11111111101010001, 17'b11111111110100001, 17'b00000000000001110, 17'b00000000000010111, 17'b11111111110111000, 17'b00000000000111101, 17'b00000000000100001, 17'b11111111111011000, 17'b11111111110010100, 17'b11111111111110110, 17'b00000000000001000, 17'b11111111111010101, 17'b00000000000001110, 17'b00000000000111010, 17'b11111111111100001, 17'b00000000000000110, 17'b00000000000000000, 17'b11111111111001000, 17'b11111111110011100, 17'b00000000001101010, 17'b00000000000100000, 17'b11111111111010010, 17'b00000000000100001, 17'b11111111111110000, 17'b11111111110000110, 17'b11111111111011101, 17'b11111111111110010, 17'b11111111111101110, 17'b00000000011010100, 17'b00000000000110000, 17'b11111111111110011, 17'b11111111111111111}, 
{17'b00000000000000011, 17'b00000000010010110, 17'b11111111101101011, 17'b11111111111000100, 17'b00000000001010010, 17'b11111111111001011, 17'b00000000100110110, 17'b11111111110110110, 17'b11111111111111111, 17'b00000000001001011, 17'b00000000001000001, 17'b11111111111111111, 17'b11111111111110011, 17'b11111111110000100, 17'b00000000001001000, 17'b00000000000101000, 17'b11111111111001110, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000001000011, 17'b11111111110001010, 17'b00000000001100100, 17'b00000000010011100, 17'b11111111111101001, 17'b11111111111111111, 17'b11111111111111011, 17'b11111111111111111, 17'b00000000010111100, 17'b00000000000000001, 17'b11111111110111010, 17'b00000000000000000, 17'b00000000001100010, 17'b11111111100110000, 17'b11111111101110101, 17'b00000000000110010, 17'b00000000000100011, 17'b11111111101101101, 17'b11111111111001111, 17'b11111111111001001, 17'b00000000001100110, 17'b00000000001100100, 17'b00000000000000000, 17'b11111111110111010, 17'b00000000000000000, 17'b00000000001100101, 17'b11111111111110000, 17'b11111111111111111, 17'b00000000000000010, 17'b00000000000111110, 17'b11111111111110001, 17'b11111111111001110, 17'b00000000001011000, 17'b11111111111001000, 17'b00000000001000111, 17'b00000000010010101, 17'b00000000000001010, 17'b00000000001000011, 17'b11111111110011001, 17'b11111111110100010, 17'b00000000011010100, 17'b11111111111011111, 17'b00000000000001011, 17'b11111111111101000}, 
{17'b00000000000000100, 17'b11111111110001100, 17'b00000000001011110, 17'b11111111110110111, 17'b11111111111111111, 17'b00000000000110110, 17'b11111111101101011, 17'b00000000000110001, 17'b00000000001111101, 17'b00000000000100111, 17'b00000000001011100, 17'b00000000001010010, 17'b11111111110110001, 17'b11111111111101100, 17'b11111111111110010, 17'b00000000000000000, 17'b11111111100001010, 17'b00000000001010010, 17'b11111111111110110, 17'b00000000000000111, 17'b11111111110100101, 17'b00000000000010001, 17'b00000000000100111, 17'b11111111111111111, 17'b11111111110001010, 17'b11111111111110011, 17'b11111111111101011, 17'b00000000100111111, 17'b11111111101010110, 17'b00000000000010001, 17'b00000000000011000, 17'b11111111111110001, 17'b11111111111000111, 17'b00000000000011101, 17'b11111111111101011, 17'b11111111111011101, 17'b11111111111010010, 17'b11111111111001010, 17'b11111111111111010, 17'b11111111110110011, 17'b00000000001010010, 17'b00000000000011111, 17'b00000000001111111, 17'b00000000000010110, 17'b00000000000001001, 17'b11111111110110101, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000000110001, 17'b00000000000101101, 17'b00000000001001011, 17'b11111111111111110, 17'b11111111110110100, 17'b00000000000000010, 17'b00000000000000000, 17'b00000000001010010, 17'b11111111111001100, 17'b11111111101110011, 17'b00000000010001111, 17'b11111111110110100, 17'b00000000100101001, 17'b11111111111111010, 17'b11111111110100101}, 
{17'b11111111101101100, 17'b11111111111111111, 17'b11111111110010111, 17'b00000000000111010, 17'b00000000001000011, 17'b11111111111100101, 17'b00000000010000100, 17'b11111111111010100, 17'b11111111110000101, 17'b11111111110100010, 17'b11111111110111111, 17'b11111111110000110, 17'b11111111111000101, 17'b00000000000110010, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000011010111, 17'b11111111111110100, 17'b11111111111111111, 17'b00000000001101001, 17'b00000000001001010, 17'b11111111101101011, 17'b11111111110011110, 17'b00000000000110000, 17'b11111111110010001, 17'b11111111111111010, 17'b11111111110111101, 17'b11111111110101010, 17'b11111111110010000, 17'b00000000001001101, 17'b00000000000111010, 17'b11111111111011000, 17'b11111111111101101, 17'b11111111100000110, 17'b11111111111010010, 17'b00000000000001100, 17'b11111111111011110, 17'b11111111110110100, 17'b11111111111111111, 17'b00000000000011110, 17'b11111111111100001, 17'b11111111111111111, 17'b11111111111110111, 17'b11111111101010101, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000001010111, 17'b11111111111100000, 17'b00000000001101100, 17'b11111111111001111, 17'b00000000001001001, 17'b11111111111111111, 17'b00000000000111001, 17'b11111111110011011, 17'b11111111111111111, 17'b00000000010000011, 17'b00000000001010000, 17'b00000000001001010, 17'b00000000000000110, 17'b11111111110011001, 17'b11111111110110011, 17'b11111111101010000, 17'b11111111111111111, 17'b00000000000011011}, 
{17'b00000000001001110, 17'b00000000000000000, 17'b00000000000100001, 17'b11111111111111111, 17'b00000000000100111, 17'b11111111111011101, 17'b00000000000111100, 17'b00000000000001010, 17'b00000000000100010, 17'b00000000001010111, 17'b11111111110111100, 17'b11111111111111010, 17'b11111111111111101, 17'b11111111111111101, 17'b11111111101010111, 17'b11111111110110011, 17'b00000000010100001, 17'b11111111111111000, 17'b11111111111110010, 17'b00000000000000000, 17'b11111111110011110, 17'b00000000000000010, 17'b00000000001000000, 17'b00000000000001001, 17'b00000000000001001, 17'b00000000001010110, 17'b00000000000000000, 17'b00000000000001001, 17'b00000000000000000, 17'b11111111111110011, 17'b11111111111001100, 17'b11111111101010101, 17'b00000000001000011, 17'b00000000001010111, 17'b11111111111111000, 17'b11111111111000011, 17'b00000000000000000, 17'b11111111101011000, 17'b11111111111110100, 17'b11111111111111111, 17'b00000000000110010, 17'b11111111111011110, 17'b11111111111111111, 17'b00000000011011000, 17'b00000000001110010, 17'b11111111111111110, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111000010, 17'b00000000000100101, 17'b00000000000100100, 17'b00000000000101100, 17'b00000000000101000, 17'b00000000001100011, 17'b00000000001011001, 17'b00000000010101000, 17'b11111111111011100, 17'b00000000001100100, 17'b00000000000100111, 17'b11111111110101100, 17'b00000000000011100, 17'b11111111110011100, 17'b11111111110001111, 17'b11111111110000000}, 
{17'b00000000000000000, 17'b00000000000111010, 17'b11111111111001110, 17'b00000000000000000, 17'b11111111111110011, 17'b11111111111110111, 17'b11111111101010110, 17'b11111111111111111, 17'b00000000001000000, 17'b00000000000111111, 17'b00000000000111100, 17'b11111111110011010, 17'b11111111111101001, 17'b00000000001001000, 17'b11111111111111111, 17'b00000000000000001, 17'b11111111100101000, 17'b11111111111111111, 17'b00000000001011111, 17'b00000000000010010, 17'b00000000000111100, 17'b11111111111100010, 17'b00000000000111111, 17'b00000000001100111, 17'b11111111110100101, 17'b11111111110111000, 17'b11111111111111110, 17'b11111111111101011, 17'b00000000000010001, 17'b00000000000000000, 17'b11111111111111111, 17'b00000000001010000, 17'b11111111101000000, 17'b00000000001011100, 17'b00000000010000000, 17'b00000000000011101, 17'b00000000000011100, 17'b11111111111100100, 17'b00000000000011101, 17'b11111111111100100, 17'b11111111110111111, 17'b11111111111110011, 17'b00000000000101010, 17'b00000000010110011, 17'b11111111100100111, 17'b11111111110001101, 17'b00000000000110001, 17'b11111111111100110, 17'b00000000001110011, 17'b11111111111000011, 17'b11111111110101011, 17'b11111111110111000, 17'b11111111111111111, 17'b00000000000011110, 17'b11111111111010111, 17'b11111111100101001, 17'b11111111111011011, 17'b11111111111111101, 17'b00000000000001011, 17'b11111111101100011, 17'b00000000100011110, 17'b11111111101110100, 17'b00000000010001010, 17'b00000000000100111}, 
{17'b00000000000010100, 17'b11111111111001110, 17'b00000000010100000, 17'b11111111110110010, 17'b11111111110001001, 17'b00000000000010111, 17'b00000000001001111, 17'b00000000001001100, 17'b11111111111010010, 17'b11111111111010110, 17'b00000000000001101, 17'b00000000000111010, 17'b00000000000111100, 17'b00000000000001100, 17'b11111111111001011, 17'b00000000000100000, 17'b00000000001111000, 17'b11111111111111101, 17'b11111111110111000, 17'b00000000000000000, 17'b00000000000010011, 17'b00000000000000101, 17'b11111111110110100, 17'b00000000000011100, 17'b00000000011001001, 17'b00000000000000010, 17'b00000000000101110, 17'b11111111100110100, 17'b11111111111101101, 17'b00000000000000010, 17'b11111111111001101, 17'b11111111110110000, 17'b00000000001110101, 17'b11111111111111001, 17'b11111111111110110, 17'b11111111110110001, 17'b00000000000100011, 17'b00000000001001010, 17'b11111111111111101, 17'b11111111111110100, 17'b11111111111010000, 17'b00000000000111010, 17'b00000000000000000, 17'b11111111101010000, 17'b00000000001001111, 17'b00000000001100110, 17'b11111111111111111, 17'b00000000000000110, 17'b11111111110010000, 17'b11111111111101100, 17'b11111111111111111, 17'b11111111110101110, 17'b00000000000000000, 17'b11111111111010011, 17'b00000000000001110, 17'b11111111100101110, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000001000110, 17'b00000000010010000, 17'b11111111101001110, 17'b00000000010000101, 17'b00000000000001001, 17'b11111111111101100}, 
{17'b00000000001001001, 17'b00000000100111101, 17'b00000000001111110, 17'b00000000001001001, 17'b11111111110000101, 17'b11111111110101110, 17'b11111110101100110, 17'b11111111110001011, 17'b00000000001100111, 17'b11111111111111111, 17'b00000000001001011, 17'b00000000011011100, 17'b00000000000010001, 17'b00000000000000001, 17'b11111111111111011, 17'b00000000000000000, 17'b11111111111001111, 17'b11111111111001100, 17'b00000000000111010, 17'b11111111101111111, 17'b11111111101010101, 17'b11111111111100101, 17'b11111111101101010, 17'b00000000000000111, 17'b11111110110111001, 17'b00000000011010000, 17'b00000000011111101, 17'b00000000010011010, 17'b11111111001000001, 17'b11111111110101111, 17'b11111111101001111, 17'b11111111100101000, 17'b11111110101111001, 17'b00000000010101101, 17'b11111111111110100, 17'b00000000001010001, 17'b00000000000000110, 17'b11111111010010001, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000000001000, 17'b00000000100000100, 17'b11111111111001011, 17'b11111111101011010, 17'b00000000011100101, 17'b11111111110001110, 17'b11111111110101100, 17'b11111111110011011, 17'b00000000001111010, 17'b00000000010001000, 17'b11111111111101110, 17'b11111111110100110, 17'b11111111111111111, 17'b11111111111100011, 17'b00000000000000000, 17'b11111111110011111, 17'b00000000010011011, 17'b00000000100010101, 17'b00000000010110110, 17'b11111111100010111, 17'b11111110001001100, 17'b00000000011100010, 17'b00000000000010111, 17'b00000000001010001}, 
{17'b11111111111000010, 17'b00000000001010110, 17'b00000000001010001, 17'b11111111111111111, 17'b11111111110100000, 17'b11111111111101001, 17'b11111111110011101, 17'b11111111111110001, 17'b00000000000100110, 17'b11111111111101100, 17'b11111111111111000, 17'b11111111111110101, 17'b11111111111111111, 17'b11111111111010001, 17'b11111111111111001, 17'b11111111111100110, 17'b00000000001010000, 17'b11111111111111111, 17'b11111111101011011, 17'b00000000001110111, 17'b00000000010011000, 17'b00000000001101010, 17'b11111111110101110, 17'b11111111111011100, 17'b11111111110100111, 17'b11111111110110101, 17'b00000000000111010, 17'b00000000000111011, 17'b00000000000111001, 17'b00000000001011100, 17'b00000000000001000, 17'b00000000001100010, 17'b11111111111110101, 17'b00000000000000001, 17'b00000000001001101, 17'b00000000000100001, 17'b11111111111101111, 17'b11111111111111101, 17'b00000000000000000, 17'b11111111110110101, 17'b11111111111000110, 17'b11111111111100011, 17'b11111111110100100, 17'b00000000001110011, 17'b00000000000000000, 17'b11111111111111110, 17'b11111111111101010, 17'b11111111111011010, 17'b11111111100110001, 17'b11111111111110110, 17'b11111111111000110, 17'b11111111111011011, 17'b11111111111100110, 17'b00000000001000011, 17'b00000000010101110, 17'b00000000000101111, 17'b11111111111111100, 17'b11111111110101000, 17'b11111111111111000, 17'b00000000000000000, 17'b00000000001010011, 17'b11111111111111010, 17'b00000000000001011, 17'b00000000000000000}
};

localparam logic signed [16:0] bias [64] = '{
17'b11111111111110110,  // -0.037350185215473175
17'b00000000001000110,  // 0.27355897426605225
17'b11111111111100000,  // -0.12378914654254913
17'b11111111111101111,  // -0.064457006752491
17'b00000000000001101,  // 0.05452875792980194
17'b00000000000011101,  // 0.11671770364046097
17'b00000000000100010,  // 0.13640816509723663
17'b00000000000010011,  // 0.07482525706291199
17'b00000000000001011,  // 0.04674031585454941
17'b11111111111001100,  // -0.20146161317825317
17'b11111111111100110,  // -0.09910125285387039
17'b00000000000100110,  // 0.15104414522647858
17'b11111111111100101,  // -0.10221704095602036
17'b11111111111011010,  // -0.1461549550294876
17'b11111111111101001,  // -0.08641516417264938
17'b00000000000101010,  // 0.16613510251045227
17'b11111111111101010,  // -0.0836295336484909
17'b11111111111110001,  // -0.05756539851427078
17'b11111111111110111,  // -0.03229188174009323
17'b11111111111111000,  // -0.028388574719429016
17'b00000000000100000,  // 0.1260243058204651
17'b11111111111110110,  // -0.037064336240291595
17'b00000000000110001,  // 0.19336333870887756
17'b00000000000000101,  // 0.02124214917421341
17'b00000000001111111,  // 0.4985624849796295
17'b00000000000000100,  // 0.0158411655575037
17'b11111111111101010,  // -0.08296407759189606
17'b00000000000011100,  // 0.11056788265705109
17'b00000000000000011,  // 0.01173810102045536
17'b11111111111100100,  // -0.10843746364116669
17'b00000000001000110,  // 0.27439257502555847
17'b00000000000010111,  // 0.09199801832437515
17'b00000000001000110,  // 0.27419957518577576
17'b00000000001000101,  // 0.27063727378845215
17'b11111111111000000,  // -0.24828937649726868
17'b00000000000010100,  // 0.07818280160427094
17'b11111111111111110,  // -0.005749030504375696
17'b00000000000011011,  // 0.10850494354963303
17'b00000000000100010,  // 0.13591453433036804
17'b11111111111100001,  // -0.12088628858327866
17'b11111111111110001,  // -0.05666546896100044
17'b00000000000010111,  // 0.09311636537313461
17'b00000000000001110,  // 0.05477767437696457
17'b00000000000000111,  // 0.029585206881165504
17'b11111111110110000,  // -0.31209176778793335
17'b11111111111101010,  // -0.08465463668107986
17'b11111111111010101,  // -0.16775836050510406
17'b00000000000100101,  // 0.14762157201766968
17'b11111111111000011,  // -0.23618532717227936
17'b00000000000010000,  // 0.06535740196704865
17'b11111111111011111,  // -0.12853026390075684
17'b11111111111011100,  // -0.13802281022071838
17'b11111111111011001,  // -0.15156887471675873
17'b00000000000010100,  // 0.07979883998632431
17'b00000000000101110,  // 0.18141601979732513
17'b11111111111110010,  // -0.054039113223552704
17'b11111111111111101,  // -0.010052933357656002
17'b00000000000010000,  // 0.06611225008964539
17'b00000000000001100,  // 0.05053366720676422
17'b00000000000000110,  // 0.026860840618610382
17'b00000000000001000,  // 0.03283466026186943
17'b00000000000100111,  // 0.15558314323425293
17'b11111111110110110,  // -0.2863388657569885
17'b11111111111101001   // -0.08769102394580841
};
endpackage