// Width: 16
// NFRAC: 6
package dense_4_16_6;

localparam logic signed [15:0] weights [32][5] = '{ 
{16'b1111111111111111, 16'b0000000000010100, 16'b1111111111101100, 16'b0000000000000100, 16'b1111111111111001}, 
{16'b1111111111011100, 16'b1111111111111100, 16'b0000000000011101, 16'b1111111111111111, 16'b0000000000000001}, 
{16'b0000000000010111, 16'b0000000000001101, 16'b1111111111111110, 16'b1111111111100110, 16'b1111111111110010}, 
{16'b1111111111100111, 16'b1111111111101000, 16'b1111111111111000, 16'b0000000000010011, 16'b0000000000001111}, 
{16'b0000000000000111, 16'b0000000000001000, 16'b0000000000001010, 16'b1111111111111110, 16'b1111111110111111}, 
{16'b0000000000010100, 16'b1111111111100110, 16'b0000000000001011, 16'b1111111111110101, 16'b1111111111110101}, 
{16'b1111111111100110, 16'b0000000000000010, 16'b1111111111111111, 16'b0000000000001011, 16'b0000000000000100}, 
{16'b1111111111111111, 16'b0000000000010010, 16'b1111111111100110, 16'b0000000000001010, 16'b0000000000001000}, 
{16'b0000000000001010, 16'b1111111111110101, 16'b0000000000000000, 16'b1111111111100010, 16'b1111111111110000}, 
{16'b1111111111111111, 16'b1111111111101110, 16'b0000000000001011, 16'b0000000000011011, 16'b0000000000000000}, 
{16'b1111111111110111, 16'b1111111111110110, 16'b0000000000000000, 16'b0000000000100101, 16'b1111111111101110}, 
{16'b0000000000001010, 16'b0000000000001110, 16'b1111111111101010, 16'b1111111111111110, 16'b0000000000000111}, 
{16'b0000000000000000, 16'b0000000000001010, 16'b0000000000000000, 16'b1111111111110010, 16'b1111111111011000}, 
{16'b0000000000001011, 16'b0000000000000100, 16'b0000000000011010, 16'b1111111111111011, 16'b1111111111100100}, 
{16'b0000000000000101, 16'b1111111111111100, 16'b1111111111101000, 16'b1111111111111101, 16'b0000000000100010}, 
{16'b1111111111100001, 16'b1111111111110000, 16'b1111111111110001, 16'b0000000000011001, 16'b0000000000000010}, 
{16'b0000000000010110, 16'b1111111111110101, 16'b1111111111110111, 16'b1111111111110001, 16'b1111111111111100}, 
{16'b0000000000001100, 16'b1111111111111101, 16'b1111111111100101, 16'b1111111111111110, 16'b0000000000000100}, 
{16'b0000000000010000, 16'b0000000000000010, 16'b1111111111110010, 16'b0000000000000000, 16'b1111111111100111}, 
{16'b0000000000001110, 16'b1111111111111010, 16'b1111111111110010, 16'b0000000000001101, 16'b0000000000000110}, 
{16'b0000000000000100, 16'b1111111111111110, 16'b0000000000010011, 16'b1111111111100100, 16'b1111111111111110}, 
{16'b0000000000000000, 16'b0000000000000111, 16'b0000000000011111, 16'b1111111111011110, 16'b1111111111011000}, 
{16'b1111111111111001, 16'b0000000000000111, 16'b0000000000001011, 16'b1111111111101001, 16'b0000000000100001}, 
{16'b1111111111111111, 16'b0000000000001010, 16'b0000000000010010, 16'b0000000000000010, 16'b1111111111011011}, 
{16'b1111111111110101, 16'b0000000000010111, 16'b1111111111110001, 16'b0000000000000000, 16'b0000000000011000}, 
{16'b0000000000000001, 16'b0000000000010001, 16'b0000000000000001, 16'b1111111111010000, 16'b0000000000100011}, 
{16'b1111111111100010, 16'b1111111111110000, 16'b0000000000001101, 16'b0000000000001111, 16'b0000000000001100}, 
{16'b0000000000000000, 16'b0000000000001111, 16'b1111111111111101, 16'b1111111111110110, 16'b0000000000000010}, 
{16'b1111111111111001, 16'b0000000000001111, 16'b1111111111011111, 16'b0000000000001000, 16'b1111111111110101}, 
{16'b1111111111111110, 16'b0000000000001001, 16'b1111111111110101, 16'b1111111111100110, 16'b0000000000100101}, 
{16'b0000000000011100, 16'b0000000000000100, 16'b0000000000010100, 16'b1111111111011010, 16'b1111111111101011}, 
{16'b1111111111111100, 16'b1111111111100111, 16'b0000000000010111, 16'b0000000000000100, 16'b0000000000001000}
};

localparam logic signed [15:0] bias [5] = '{
16'b1111111111111100,  // -0.06223141402006149
16'b1111111111111011,  // -0.06270556896924973
16'b1111111111111011,  // -0.07014333456754684
16'b0000000000000101,  // 0.0820775106549263
16'b0000000000001101   // 0.2155742198228836
};
endpackage