// Width: 15
// NFRAC: 7
package dense_4_15_7;

localparam logic signed [14:0] weights [32][5] = '{ 
{15'b111111111111110, 15'b000000000101000, 15'b111111111011001, 15'b000000000001000, 15'b111111111110010}, 
{15'b111111110111000, 15'b111111111111000, 15'b000000000111010, 15'b111111111111110, 15'b000000000000010}, 
{15'b000000000101111, 15'b000000000011011, 15'b111111111111100, 15'b111111111001100, 15'b111111111100101}, 
{15'b111111111001111, 15'b111111111010000, 15'b111111111110001, 15'b000000000100111, 15'b000000000011110}, 
{15'b000000000001111, 15'b000000000010000, 15'b000000000010100, 15'b111111111111101, 15'b111111101111110}, 
{15'b000000000101001, 15'b111111111001101, 15'b000000000010111, 15'b111111111101011, 15'b111111111101010}, 
{15'b111111111001100, 15'b000000000000100, 15'b111111111111111, 15'b000000000010110, 15'b000000000001000}, 
{15'b111111111111111, 15'b000000000100100, 15'b111111111001101, 15'b000000000010100, 15'b000000000010001}, 
{15'b000000000010100, 15'b111111111101010, 15'b000000000000000, 15'b111111111000100, 15'b111111111100000}, 
{15'b111111111111111, 15'b111111111011101, 15'b000000000010110, 15'b000000000110111, 15'b000000000000000}, 
{15'b111111111101111, 15'b111111111101101, 15'b000000000000000, 15'b000000001001010, 15'b111111111011101}, 
{15'b000000000010101, 15'b000000000011101, 15'b111111111010100, 15'b111111111111100, 15'b000000000001111}, 
{15'b000000000000000, 15'b000000000010101, 15'b000000000000001, 15'b111111111100101, 15'b111111110110000}, 
{15'b000000000010110, 15'b000000000001000, 15'b000000000110101, 15'b111111111110111, 15'b111111111001001}, 
{15'b000000000001011, 15'b111111111111001, 15'b111111111010001, 15'b111111111111011, 15'b000000001000100}, 
{15'b111111111000011, 15'b111111111100000, 15'b111111111100011, 15'b000000000110011, 15'b000000000000100}, 
{15'b000000000101100, 15'b111111111101010, 15'b111111111101110, 15'b111111111100011, 15'b111111111111000}, 
{15'b000000000011000, 15'b111111111111010, 15'b111111111001011, 15'b111111111111100, 15'b000000000001001}, 
{15'b000000000100001, 15'b000000000000101, 15'b111111111100100, 15'b000000000000000, 15'b111111111001111}, 
{15'b000000000011101, 15'b111111111110100, 15'b111111111100100, 15'b000000000011010, 15'b000000000001100}, 
{15'b000000000001000, 15'b111111111111100, 15'b000000000100110, 15'b111111111001000, 15'b111111111111101}, 
{15'b000000000000000, 15'b000000000001111, 15'b000000000111110, 15'b111111110111101, 15'b111111110110000}, 
{15'b111111111110011, 15'b000000000001110, 15'b000000000010110, 15'b111111111010010, 15'b000000001000010}, 
{15'b111111111111111, 15'b000000000010101, 15'b000000000100100, 15'b000000000000100, 15'b111111110110110}, 
{15'b111111111101010, 15'b000000000101110, 15'b111111111100011, 15'b000000000000000, 15'b000000000110001}, 
{15'b000000000000011, 15'b000000000100010, 15'b000000000000011, 15'b111111110100000, 15'b000000001000110}, 
{15'b111111111000101, 15'b111111111100000, 15'b000000000011011, 15'b000000000011111, 15'b000000000011001}, 
{15'b000000000000000, 15'b000000000011110, 15'b111111111111011, 15'b111111111101100, 15'b000000000000100}, 
{15'b111111111110010, 15'b000000000011111, 15'b111111110111111, 15'b000000000010001, 15'b111111111101011}, 
{15'b111111111111101, 15'b000000000010010, 15'b111111111101010, 15'b111111111001100, 15'b000000001001011}, 
{15'b000000000111001, 15'b000000000001000, 15'b000000000101001, 15'b111111110110100, 15'b111111111010111}, 
{15'b111111111111000, 15'b111111111001110, 15'b000000000101110, 15'b000000000001001, 15'b000000000010000}
};

localparam logic signed [14:0] bias [5] = '{
15'b111111111111000,  // -0.06223141402006149
15'b111111111110111,  // -0.06270556896924973
15'b111111111110111,  // -0.07014333456754684
15'b000000000001010,  // 0.0820775106549263
15'b000000000011011   // 0.2155742198228836
};
endpackage