// Width: 23
// NFRAC: 11
package dense_2_23_11;

localparam logic signed [22:0] weights [64][32] = '{ 
{23'b00000000000001000100110, 23'b00000000000000000010000, 23'b11111111111111001111011, 23'b11111111111111111010100, 23'b00000000000001000010110, 23'b00000000000000000000000, 23'b11111111111111011011000, 23'b11111111111111111111111, 23'b11111111111110111001111, 23'b00000000000000010100011, 23'b00000000000000000000000, 23'b11111111111111111110100, 23'b11111111111111111111111, 23'b11111111111111001100110, 23'b11111111111111110011000, 23'b11111111111110111100111, 23'b00000000000000000000000, 23'b11111111111111111100101, 23'b11111111111111001111001, 23'b11111111111111010111011, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b11111111111111111101111, 23'b11111111111111111111010, 23'b00000000000000000000000, 23'b00000000000000011001101, 23'b00000000000001100010110, 23'b00000000000000101100110, 23'b11111111111111111111111, 23'b00000000000000001100111, 23'b11111111111110010111001, 23'b00000000000000000000000}, 
{23'b11111111111111100110010, 23'b11111111111111011000010, 23'b11111111111111011100100, 23'b11111111111111110001110, 23'b11111111111111111110100, 23'b00000000000000001011000, 23'b11111111111111000110110, 23'b00000000000000000001010, 23'b00000000000000000001001, 23'b11111111111111101111111, 23'b00000000000000100111111, 23'b11111111111111110100111, 23'b11111111111111110000111, 23'b11111111111111001000011, 23'b00000000000000000001111, 23'b11111111111111110011101, 23'b00000000000000000011001, 23'b11111111111111001110001, 23'b00000000000000101011111, 23'b00000000000000111010110, 23'b11111111111111110111111, 23'b11111111111111111110100, 23'b11111111111111111111111, 23'b00000000000000000110000, 23'b11111111111111101101110, 23'b00000000000001000110011, 23'b00000000000000111111011, 23'b00000000000000000010001, 23'b00000000000000000111010, 23'b11111111111110000011011, 23'b00000000000000000001111, 23'b00000000000000000000000}, 
{23'b00000000000000010010100, 23'b11111111111111100010101, 23'b11111111111111011110110, 23'b11111111111111110101010, 23'b11111111111111101100001, 23'b11111111111111101010001, 23'b11111111111111010000101, 23'b00000000000000000001001, 23'b11111111111111011101011, 23'b00000000000000000010010, 23'b00000000000000000000100, 23'b11111111111111101011010, 23'b00000000000000010111001, 23'b11111111111111101111011, 23'b11111111111111111111101, 23'b11111111111111110110100, 23'b00000000000000000001010, 23'b00000000000000011000011, 23'b00000000000000001111000, 23'b00000000000000111010110, 23'b00000000000000001010100, 23'b11111111111111101010011, 23'b00000000000000000000000, 23'b00000000000000001000111, 23'b11111111111111111011010, 23'b00000000000000110101100, 23'b00000000000000100110001, 23'b00000000000000011000110, 23'b11111111111111111111111, 23'b11111111111111011001000, 23'b11111111111111111100100, 23'b00000000000000011001011}, 
{23'b00000000000000100011010, 23'b00000000000000000100111, 23'b00000000000000001101100, 23'b11111111111111111101100, 23'b11111111111101111101101, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b00000000000000111001111, 23'b00000000000000111110000, 23'b11111111111111111100100, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b00000000000000000001010, 23'b11111111111111111011010, 23'b00000000000000110110111, 23'b00000000000000000000000, 23'b11111111111111111001101, 23'b11111111111111111111111, 23'b11111111111111010010111, 23'b11111111111111110000010, 23'b00000000000000001100101, 23'b11111111111111101111110, 23'b11111111111111111111111, 23'b00000000000000000000111, 23'b11111111111111110011000, 23'b00000000000000010010101, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b11111111111111001000111, 23'b00000000000001001111011}, 
{23'b11111111111101010001010, 23'b11111111111111111001101, 23'b11111111111111111110111, 23'b00000000000000000001010, 23'b11111111111111111001010, 23'b00000000000000000001101, 23'b11111111111111110011011, 23'b11111111111111011001101, 23'b00000000000000001101111, 23'b11111111111111111010110, 23'b11111111111111111100100, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b00000000000000110101110, 23'b00000000000000000000000, 23'b00000000000001010100001, 23'b11111111111111111111111, 23'b00000000000000110111110, 23'b11111111111110011001100, 23'b00000000000000000000000, 23'b11111111111111100011011, 23'b00000000000000101011001, 23'b00000000000001000010000, 23'b00000000000000000000000, 23'b00000000000000001011100, 23'b00000000000000101001101, 23'b00000000000000111101000, 23'b00000000000000000100011, 23'b11111111111111111110110, 23'b11111111111111111111111, 23'b11111111111111111100011, 23'b00000000000000111001111}, 
{23'b00000000000000001110110, 23'b11111111111111111111111, 23'b00000000000000100110001, 23'b11111111111101011001111, 23'b11111111111010011111011, 23'b11111111111110100110010, 23'b00000000000001011010101, 23'b11111111111101100000101, 23'b11111111111111111111111, 23'b11111111111101010010100, 23'b11111111111101111111101, 23'b11111111111110101000101, 23'b00000000000001011010011, 23'b11111111111111111111111, 23'b11111111111111111100001, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b11111111111111011110001, 23'b11111111111111111111111, 23'b11111111111110000010110, 23'b00000000000000000000000, 23'b00000000000000101111100, 23'b11111111111111111111111, 23'b00000000000000000101101, 23'b00000000000001000100100, 23'b00000000000000001101000, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b00000000000000110100101, 23'b11111111111111110111010, 23'b00000000000000110011010}, 
{23'b11111111111111110110110, 23'b11111111111111010111101, 23'b11111111111111000010001, 23'b11111111111111110011111, 23'b11111111111110110110001, 23'b00000000000000010000111, 23'b11111111111111010001111, 23'b11111111111111011011101, 23'b11111111111110010101110, 23'b00000000000000001100011, 23'b11111111111111111110101, 23'b11111111111111010111010, 23'b00000000000000011110011, 23'b11111111111111111101011, 23'b11111111111111110101011, 23'b11111111111101110010010, 23'b11111111111111111111111, 23'b00000000000000010101100, 23'b00000000000000110001000, 23'b11111111111111010110011, 23'b11111111111111011001100, 23'b11111111111111101111111, 23'b11111111111111111111101, 23'b00000000000000000111000, 23'b11111111111111110100010, 23'b11111111111101011010000, 23'b11111111111110111100001, 23'b11111111111111110100011, 23'b00000000000000000001011, 23'b11111111111111111010100, 23'b00000000000000000111110, 23'b11111111111111111111110}, 
{23'b11111111111111011000101, 23'b11111111111111101000110, 23'b11111111111111101011101, 23'b11111111111111000011010, 23'b11111111111111100010010, 23'b11111111111111111111111, 23'b00000000000000011010101, 23'b11111111111111101011110, 23'b00000000000000110011010, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b00000000000000111000000, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b11111111111111101101111, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b11111111111111111111110, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b00000000000000001011010, 23'b11111111111111010001111, 23'b00000000000000000011100, 23'b11111111111111111111111, 23'b11111111111111101101100, 23'b11111111111111111111110, 23'b00000000000000000000000, 23'b11111111111111111111111}, 
{23'b11111111111110000101110, 23'b11111111111111110001011, 23'b11111111111110011110101, 23'b00000000000000011111010, 23'b00000000000001111100101, 23'b11111111111111111111111, 23'b11111111111111111000100, 23'b00000000000000111101001, 23'b11111111111110001111101, 23'b11111111111111110100000, 23'b00000000000000000000000, 23'b11111111111111001100011, 23'b11111111111111111111111, 23'b00000000000000010011011, 23'b11111111111111001111001, 23'b00000000000011000001000, 23'b11111111111111111101110, 23'b00000000000000001011111, 23'b00000000000000110101001, 23'b00000000000000111110101, 23'b00000000000000000000000, 23'b11111111111110101010000, 23'b00000000000000000000000, 23'b00000000000001101001010, 23'b11111111111111010001100, 23'b00000000000010110010100, 23'b11111111111111011001110, 23'b11111111111111001011110, 23'b11111111111110000111001, 23'b11111111111110001001001, 23'b00000000000000000000000, 23'b00000000000000001101101}, 
{23'b00000000000000000000000, 23'b11111111111111111100000, 23'b11111111111111101101000, 23'b00000000000000000000000, 23'b00000000000001001110111, 23'b11111111111111111010110, 23'b11111111111111101111101, 23'b00000000000000010111100, 23'b00000000000000011001111, 23'b00000000000000000000111, 23'b11111111111111111101110, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b11111111111111100010111, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b11111111111111111110101, 23'b00000000000000000000100, 23'b00000000000000010101101, 23'b00000000000000000100111, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b00000000000000000001110, 23'b00000000000000001001110, 23'b11111111111111011110001, 23'b00000000000000010001011, 23'b00000000000000111111101, 23'b11111111111111111111111, 23'b00000000000000000001100, 23'b00000000000000001100101, 23'b00000000000000010001110}, 
{23'b00000000000000011000101, 23'b00000000000000000000000, 23'b11111111111111100101100, 23'b11111111111110111111110, 23'b11111111111100110100101, 23'b00000000000000100010000, 23'b00000000000000000000000, 23'b11111111111100101100001, 23'b00000000000000001001010, 23'b11111111111111111111111, 23'b00000000000000000000111, 23'b11111111111111111111100, 23'b00000000000000000010101, 23'b00000000000000000000000, 23'b11111111111111111011001, 23'b11111111111110011110010, 23'b11111111111111111111111, 23'b00000000000000111000010, 23'b00000000000000100000010, 23'b00000000000000110000111, 23'b11111111111110001111011, 23'b11111111111110100100111, 23'b00000000000000011110101, 23'b11111111111111110111000, 23'b11111111111111110100001, 23'b00000000000001011011110, 23'b11111111111111100111010, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b00000000000000110110000, 23'b11111111111111111111111, 23'b00000000000000000001100}, 
{23'b11111111111111001101011, 23'b11111111111110000001110, 23'b00000000000000000000000, 23'b11111111111111111111011, 23'b00000000000001010101000, 23'b11111111111110111011000, 23'b11111111111111000111010, 23'b00000000000000011101101, 23'b11111111111111111111110, 23'b00000000000000100110000, 23'b00000000000000010010111, 23'b11111111111111101100101, 23'b00000000000000000000000, 23'b00000000000000000011100, 23'b11111111111111111010100, 23'b11111111111110111111001, 23'b00000000000000101100111, 23'b00000000000000000111010, 23'b00000000000001001100000, 23'b00000000000000010110001, 23'b00000000000000000000000, 23'b11111111111111110110010, 23'b00000000000000100000010, 23'b11111111111111101001111, 23'b11111111111110110001001, 23'b11111111111111111110010, 23'b00000000000000101111010, 23'b11111111111111111111111, 23'b00000000000000000010001, 23'b11111111111111100111110, 23'b00000000000000100011001, 23'b00000000000001000110101}, 
{23'b00000000000000000011111, 23'b00000000000000000000000, 23'b00000000000000111000001, 23'b00000000000000000010001, 23'b11111111111111110101100, 23'b00000000000000101110001, 23'b00000000000000010111100, 23'b11111111111111111111111, 23'b00000000000000000000001, 23'b11111111111111011100000, 23'b11111111111111110010000, 23'b11111111111111010101001, 23'b11111111111111111111111, 23'b00000000000000001100111, 23'b11111111111111101110010, 23'b00000000000011010111110, 23'b00000000000000000000000, 23'b11111111111111100111111, 23'b11111111111111001111101, 23'b11111111111111111100100, 23'b00000000000000110010110, 23'b00000000000000100000110, 23'b00000000000000000000000, 23'b11111111111111111111010, 23'b00000000000000111000001, 23'b00000000000001000100101, 23'b00000000000001111110110, 23'b00000000000000000010101, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b11111111111111111100111, 23'b11111111111111101101101}, 
{23'b11111111111111011000000, 23'b00000000000000001100011, 23'b00000000000000001010000, 23'b11111111111111000000101, 23'b11111111111110111011000, 23'b00000000000001111000000, 23'b00000000000000001100100, 23'b00000000000000000000000, 23'b11111111111111010110110, 23'b11111111111111101001011, 23'b00000000000000100001001, 23'b00000000000000010010001, 23'b00000000000000000000001, 23'b11111111111111101011111, 23'b00000000000001001001001, 23'b11111111111111111111111, 23'b11111111111111111100100, 23'b00000000000000000000000, 23'b00000000000000000011010, 23'b11111111111111110100000, 23'b00000000000000010100000, 23'b00000000000000000100000, 23'b00000000000000011101001, 23'b11111111111111111111111, 23'b00000000000000000000110, 23'b00000000000010101000011, 23'b11111111111111110001100, 23'b11111111111111111010000, 23'b11111111111111111111111, 23'b11111111111111100100000, 23'b11111111111111110101101, 23'b00000000000000101101000}, 
{23'b00000000000000001111000, 23'b00000000000000010010111, 23'b00000000000001010011100, 23'b11111111111111110101110, 23'b00000000000000011001110, 23'b00000000000001011001110, 23'b00000000000000000000001, 23'b11111111111111111000011, 23'b00000000000000011110001, 23'b11111111111111100010110, 23'b11111111111111111111111, 23'b11111111111111100001011, 23'b00000000000000000000000, 23'b00000000000001100100101, 23'b11111111111111111011011, 23'b00000000000000000000011, 23'b00000000000000111100011, 23'b00000000000000000000001, 23'b00000000000000000000110, 23'b11111111111110101111111, 23'b11111111111111000001001, 23'b11111111111111110110110, 23'b11111111111111111111111, 23'b11111111111111011010101, 23'b11111111111111110110110, 23'b11111111111111101010111, 23'b11111111111111001101101, 23'b11111111111111001001100, 23'b00000000000000000111101, 23'b00000000000000011100100, 23'b11111111111110011010010, 23'b00000000000000000000110}, 
{23'b11111111111110110011100, 23'b00000000000000000000000, 23'b11111111111111111100001, 23'b11111111111111110011010, 23'b11111111111111111111111, 23'b00000000000000100010001, 23'b11111111111111101100001, 23'b00000000000001000101011, 23'b11111111111110100011000, 23'b11111111111111111111110, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b11111111111111111111000, 23'b11111111111111101000110, 23'b00000000000000010100010, 23'b00000000000000101110111, 23'b11111111111111111101100, 23'b11111111111110111111101, 23'b11111111111111110000111, 23'b00000000000000011100101, 23'b00000000000000010000001, 23'b00000000000000000000000, 23'b00000000000000000000110, 23'b00000000000000010100111, 23'b11111111111111000010101, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b00000000000000000000110, 23'b00000000000000000000001, 23'b11111111111111011111110}, 
{23'b11111111111110101001111, 23'b11111111111111111110100, 23'b11111111111111111111001, 23'b11111111111111111011100, 23'b11111111111111111110110, 23'b00000000000000011011000, 23'b00000000000000000001101, 23'b00000000000000001000110, 23'b00000000000000001001110, 23'b00000000000000010000000, 23'b00000000000000010100001, 23'b00000000000000101001010, 23'b00000000000000000110110, 23'b11111111111111100111001, 23'b00000000000000000000001, 23'b00000000000001100001101, 23'b00000000000000000000000, 23'b00000000000000000000010, 23'b11111111111111111111010, 23'b00000000000000011100001, 23'b00000000000000100100011, 23'b00000000000000000111111, 23'b00000000000000001010100, 23'b11111111111111111000011, 23'b11111111111111110111110, 23'b00000000000000000110110, 23'b11111111111111101110110, 23'b11111111111111011111100, 23'b00000000000000110101101, 23'b11111111111111111000001, 23'b00000000000000001000000, 23'b11111111111111001111111}, 
{23'b00000000000000000000000, 23'b11111111111111111111111, 23'b00000000000000001001101, 23'b00000000000000000000000, 23'b00000000000011101000000, 23'b11111111111111111111110, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b00000000000000011100000, 23'b11111111111111101100110, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b00000000000000000000010, 23'b00000000000000100001000, 23'b00000000000000000000000, 23'b11111111111111011010110, 23'b11111111111111111111111, 23'b11111111111111101110110, 23'b00000000000001010011110, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b00000000000000010001011, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b00000000000000001010100}, 
{23'b11111111111111111111001, 23'b00000000000000000111011, 23'b11111111111111111111110, 23'b00000000000000001100010, 23'b11111111111111110100101, 23'b11111111111111100001011, 23'b11111111111111110000000, 23'b00000000000001000111000, 23'b00000000000000000000000, 23'b00000000000000011000110, 23'b11111111111111111101001, 23'b00000000000000010000100, 23'b11111111111111110111100, 23'b11111111111111010111101, 23'b11111111111111001111001, 23'b00000000000000000011010, 23'b11111111111111111111111, 23'b11111111111111110111000, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b11111111111111111111110, 23'b00000000000000010011011, 23'b00000000000000001001001, 23'b11111111111111011111110, 23'b00000000000000011100100, 23'b11111111111111010101111, 23'b00000000000000000000100, 23'b00000000000000000000000, 23'b11111111111111010101000, 23'b00000000000000000000000, 23'b00000000000000001011101, 23'b11111111111111111000000}, 
{23'b11111111111111111101000, 23'b11111111111111100110101, 23'b00000000000000000000000, 23'b11111111111111110000101, 23'b00000000000000110111010, 23'b11111111111111111111111, 23'b11111111111111111010101, 23'b00000000000000011011010, 23'b11111111111110011011111, 23'b00000000000000000000000, 23'b11111111111111110110001, 23'b11111111111111111111011, 23'b00000000000001011001111, 23'b00000000000000111010101, 23'b11111111111111100110100, 23'b11111111111111111010101, 23'b11111111111111111111111, 23'b00000000000000000000001, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b11111111111111011101001, 23'b11111111111111100001100, 23'b00000000000000100001100, 23'b00000000000000000000000, 23'b11111111111111011100111, 23'b00000000000000000110010, 23'b11111111111111101011011, 23'b11111111111111110111011, 23'b00000000000000100010110, 23'b00000000000000000000001, 23'b11111111111111000000101}, 
{23'b00000000000010100010011, 23'b00000000000001010111100, 23'b11111111111111000000001, 23'b00000000000000000000110, 23'b11111111111110100111011, 23'b00000000000000000000000, 23'b00000000000000111001000, 23'b00000000000000000111111, 23'b00000000000000111001010, 23'b11111111111111111111111, 23'b11111111111111011000010, 23'b11111111111111101011111, 23'b00000000000000100100010, 23'b00000000000000000111000, 23'b11111111111111100110110, 23'b00000000000000100001101, 23'b00000000000010001001000, 23'b11111111111111011110101, 23'b11111111111110110100001, 23'b00000000000000000000000, 23'b11111111111111111000101, 23'b11111111111111010010110, 23'b11111111111111111100111, 23'b11111111111111111111100, 23'b00000000000000010110000, 23'b11111111111110100011101, 23'b00000000000000010110110, 23'b11111111111111111111101, 23'b00000000000000000000000, 23'b00000000000000011011111, 23'b11111111111111111000100, 23'b00000000000000001111010}, 
{23'b11111111111111101000010, 23'b11111111111111001110110, 23'b11111111111111110110101, 23'b11111111111111010101001, 23'b11111111111111111011100, 23'b00000000000000001100100, 23'b00000000000000000000000, 23'b11111111111111111101000, 23'b00000000000000001001101, 23'b11111111111111111111000, 23'b00000000000000000000000, 23'b11111111111111001000011, 23'b00000000000000011010000, 23'b00000000000000010100100, 23'b11111111111111100101110, 23'b00000000000001110001100, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b11111111111111111110111, 23'b00000000000000000000000, 23'b00000000000001010000111, 23'b11111111111110000111100, 23'b11111111111111100100010, 23'b11111111111111110001101, 23'b11111111111111111011001, 23'b00000000000000110010011, 23'b11111111111111110010100, 23'b00000000000000000100100, 23'b00000000000001111011111, 23'b11111111111101111100110, 23'b11111111111110100010000, 23'b00000000000000000101101}, 
{23'b00000000000000000100010, 23'b11111111111111110000111, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b11111111111101000111111, 23'b11111111111101100100110, 23'b00000000000000000000011, 23'b11111111111111111111111, 23'b11111111111110111100001, 23'b00000000000000000110010, 23'b00000000000000000000000, 23'b11111111111111111000111, 23'b00000000000000000000000, 23'b11111111111111110001000, 23'b11111111111111110010100, 23'b11111111111111101110010, 23'b11111111111111011010010, 23'b00000000000001001000010, 23'b00000000000000000000000, 23'b00000000000000001011110, 23'b11111111111111111111111, 23'b11111111111111101101111, 23'b00000000000000000000000, 23'b11111111111111101001110, 23'b00000000000000111000001, 23'b11111111111101100000101, 23'b00000000000000111000010, 23'b11111111111111111111111, 23'b11111111111111111110110, 23'b00000000000000110011001, 23'b11111111111111111111111, 23'b00000000000000111100011}, 
{23'b11111111111111111111111, 23'b00000000000000000001010, 23'b11111111111111110100111, 23'b00000000000000010011001, 23'b00000000000000001110001, 23'b11111111111110101000011, 23'b00000000000000000000000, 23'b00000000000000010000011, 23'b00000000000010010100011, 23'b11111111111111111101101, 23'b00000000000000000000000, 23'b00000000000000001110011, 23'b00000000000001011011111, 23'b11111111111111110111110, 23'b00000000000000000011100, 23'b00000000000000011001110, 23'b11111111111111111111111, 23'b00000000000000000111000, 23'b11111111111111111111111, 23'b00000000000000000000001, 23'b11111111111110111001111, 23'b00000000000000001001110, 23'b00000000000000010001111, 23'b00000000000000000101110, 23'b11111111111111111111111, 23'b00000000000000110111111, 23'b00000000000000000001001, 23'b00000000000000100000010, 23'b11111111111110010101000, 23'b00000000000000011010010, 23'b00000000000001100101010, 23'b00000000000000000001011}, 
{23'b11111111111110100110001, 23'b00000000000000110110000, 23'b11111111111110111101010, 23'b00000000000000011111011, 23'b11111111111111100101000, 23'b00000000000000000000000, 23'b00000000000001111111011, 23'b11111111111111000100011, 23'b11111111111110110101011, 23'b00000000000000101011110, 23'b11111111111111000110111, 23'b11111111111111111001111, 23'b11111111111111111111110, 23'b00000000000001011000000, 23'b11111111111111111111100, 23'b11111111111110110010110, 23'b11111111111111111111111, 23'b00000000000001110000110, 23'b11111111111110000111011, 23'b11111111111111111001110, 23'b00000000000001010001000, 23'b11111111111110100011001, 23'b00000000000000001101100, 23'b11111111111111111100001, 23'b00000000000001000101011, 23'b11111111111101111101110, 23'b11111111111110100011001, 23'b11111111111111001101110, 23'b11111111111111111111111, 23'b00000000000000011010100, 23'b00000000000000000110011, 23'b00000000000000101101101}, 
{23'b11111111111111101000110, 23'b00000000000000001101010, 23'b11111111111111111111111, 23'b00000000000000100110010, 23'b11111111111111110110010, 23'b00000000000000111010000, 23'b00000000000000000000100, 23'b11111111111111111101001, 23'b11111111111111111111011, 23'b00000000000000000000010, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b11111111111111111111100, 23'b00000000000010000101001, 23'b00000000000000000011001, 23'b00000000000000110000010, 23'b00000000000000000000000, 23'b11111111111111001001110, 23'b11111111111111101100011, 23'b11111111111111111111111, 23'b11111111111111111011110, 23'b00000000000000001010110, 23'b11111111111111111111111, 23'b11111111111111010000100, 23'b11111111111111111111111, 23'b00000000000001001011101, 23'b00000000000001001111011, 23'b11111111111111111111111, 23'b11111111111111111011110, 23'b00000000000000000000000, 23'b11111111111111111111110, 23'b11111111111111100111010}, 
{23'b11111111111111101011010, 23'b00000000000000000000000, 23'b00000000000001000101111, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b11111111111111100010111, 23'b00000000000000000000000, 23'b11111111111100100010111, 23'b00000000000000110111001, 23'b00000000000000000011100, 23'b00000000000000000110110, 23'b11111111111110100011111, 23'b00000000000000000000110, 23'b11111111111111011100110, 23'b11111111111111110111100, 23'b00000000000000000000000, 23'b00000000000000000101000, 23'b00000000000000000000000, 23'b00000000000000011100110, 23'b00000000000000000000000, 23'b11111111111111111101101, 23'b00000000000001010100010, 23'b00000000000001100000011, 23'b11111111111111000111011, 23'b11111111111111011011101, 23'b00000000000000111111111, 23'b11111111111110110001110, 23'b00000000000000000111100, 23'b11111111111111111111110, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b00000000000000101111001}, 
{23'b11111111111111100010111, 23'b11111111111111111111110, 23'b11111111111111000010110, 23'b11111111111111001100010, 23'b11111111111111111100011, 23'b11111111111111011101011, 23'b00000000000000000000000, 23'b00000000000000010111010, 23'b11111111111111000010101, 23'b11111111111111101010101, 23'b11111111111111110011010, 23'b00000000000000000000000, 23'b00000000000000000111001, 23'b11111111111111111101011, 23'b11111111111111110000011, 23'b00000000000000011000011, 23'b00000000000000111001000, 23'b00000000000000100001100, 23'b11111111111111011110100, 23'b00000000000000001100011, 23'b11111111111111111100111, 23'b11111111111111111000101, 23'b00000000000000000101110, 23'b00000000000000000100000, 23'b11111111111111101110001, 23'b00000000000000010110110, 23'b11111111111111101000110, 23'b00000000000000001111010, 23'b11111111111111111111111, 23'b11111111111110110100011, 23'b11111111111111111001010, 23'b00000000000000111001100}, 
{23'b11111111111111111001000, 23'b11111111111111101010110, 23'b00000000000000010011101, 23'b00000000000001000000110, 23'b00000000000000010101101, 23'b00000000000000010101000, 23'b00000000000000001011111, 23'b11111111111111001100011, 23'b11111111111111001011011, 23'b00000000000000010001100, 23'b00000000000000000011000, 23'b00000000000000001011000, 23'b00000000000000000101101, 23'b00000000000000000001011, 23'b00000000000000110100100, 23'b00000000000000000001111, 23'b11111111111111110010001, 23'b00000000000000011010011, 23'b11111111111111111000011, 23'b11111111111111110110110, 23'b00000000000000011100001, 23'b11111111111111100000010, 23'b11111111111111111001001, 23'b00000000000000100000100, 23'b00000000000000000101101, 23'b11111111111111100100101, 23'b11111111111111001101010, 23'b11111111111111111100111, 23'b11111111111110111000100, 23'b00000000000000001111011, 23'b00000000000000011010000, 23'b00000000000000000000010}, 
{23'b11111111111111111100100, 23'b11111111111111111010111, 23'b11111111111111111100111, 23'b11111111111111110111001, 23'b11111111111111011110010, 23'b11111111111111011100000, 23'b00000000000000010000001, 23'b00000000000000000010000, 23'b11111111111111010001010, 23'b00000000000000101010110, 23'b11111111111111111010101, 23'b11111111111111111111110, 23'b11111111111111100011110, 23'b00000000000000000001010, 23'b00000000000000000111100, 23'b11111111111111110010100, 23'b11111111111111111011111, 23'b11111111111111110101010, 23'b11111111111111101011011, 23'b00000000000000000000000, 23'b11111111111111011100000, 23'b00000000000000011010000, 23'b11111111111111001001110, 23'b00000000000000000001010, 23'b00000000000000001010101, 23'b00000000000000011111101, 23'b00000000000000000110110, 23'b00000000000000000001100, 23'b00000000000001001010110, 23'b00000000000000001101001, 23'b00000000000000000000000, 23'b00000000000000010101011}, 
{23'b11111111111111111011000, 23'b00000000000001000000101, 23'b11111111111111111111111, 23'b11111111111111110111100, 23'b11111111111111001001010, 23'b11111111111111101100110, 23'b00000000000001101001010, 23'b11111111111101001111100, 23'b11111111111110100110100, 23'b11111111111111001100111, 23'b11111111111111000111110, 23'b11111111111110111111000, 23'b11111111111111111111110, 23'b00000000000001111011111, 23'b11111111111111111001010, 23'b00000000000000000000000, 23'b11111111111111001001111, 23'b00000000000001110010000, 23'b11111111111110010110010, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b11111111111110101001111, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b00000000000000001110011, 23'b11111111111111110001010, 23'b11111111111111011010001, 23'b11111111111111111111111, 23'b00000000000000101100101, 23'b00000000000000000000110, 23'b11111111111111101011011, 23'b00000000000000000000001}, 
{23'b00000000000001011110001, 23'b11111111111111100011010, 23'b00000000000000100001110, 23'b11111111111111110111101, 23'b00000000000000010011100, 23'b11111111111111111111000, 23'b11111111111111111111010, 23'b11111111111111101000001, 23'b00000000000000000000000, 23'b00000000000000010111100, 23'b11111111111111111111111, 23'b11111111111111110000111, 23'b11111111111111111111111, 23'b00000000000000111010100, 23'b00000000000000000100111, 23'b00000000000000001010010, 23'b00000000000000000110001, 23'b11111111111111111001110, 23'b00000000000000000101001, 23'b00000000000000000000000, 23'b11111111111111111101101, 23'b11111111111111111111111, 23'b11111111111110110001110, 23'b11111111111111111111111, 23'b00000000000000001110110, 23'b11111111111111100010001, 23'b11111111111111011101011, 23'b11111111111111111111111, 23'b11111111111111111111110, 23'b00000000000010001110110, 23'b11111111111110110110110, 23'b11111111111111100010010}, 
{23'b11111111111111110100101, 23'b11111111111111100101100, 23'b11111111111111101111011, 23'b00000000000000001001010, 23'b00000000000000100011101, 23'b11111111111111011110110, 23'b11111111111111111111101, 23'b11111111111111000111101, 23'b00000000000000001111100, 23'b00000000000000100010110, 23'b11111111111111001001010, 23'b11111111111110111111010, 23'b00000000000000000110000, 23'b11111111111101010001000, 23'b11111111111111101100101, 23'b11111111111111100000011, 23'b11111111111111001101010, 23'b11111111111111111111111, 23'b00000000000000100010010, 23'b00000000000000000000000, 23'b11111111111111110100010, 23'b11111111111111110100100, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b11111111111111110000111, 23'b11111111111100111110111, 23'b11111111111101110001110, 23'b11111111111110111010001, 23'b00000000000000001110010, 23'b00000000000000110100110, 23'b11111111111111111111111, 23'b00000000000000111101100}, 
{23'b11111111111111101000011, 23'b11111111111111001001000, 23'b00000000000000101001111, 23'b00000000000000010011000, 23'b00000000000000001011000, 23'b11111111111111101000011, 23'b11111111111111110111101, 23'b00000000000000011001001, 23'b00000000000010001001111, 23'b11111111111111010100001, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b00000000000000011110000, 23'b11111111111111110001111, 23'b11111111111111111011011, 23'b11111111111111111011101, 23'b11111111111111100110011, 23'b11111111111111111111110, 23'b00000000000000000000000, 23'b00000000000000111010000, 23'b11111111111111011101111, 23'b11111111111111111111001, 23'b00000000000000100000111, 23'b11111111111111111101011, 23'b00000000000000000000000, 23'b00000000000010000110101, 23'b00000000000001010011000, 23'b00000000000000000000110, 23'b00000000000000000000000, 23'b11111111111110010100010, 23'b11111111111111101110100, 23'b11111111111111111111111}, 
{23'b00000000000000000011110, 23'b00000000000000001100010, 23'b11111111111111111100011, 23'b00000000000000000000000, 23'b00000000000000111011001, 23'b11111111111110000100010, 23'b00000000000000000000000, 23'b11111111111111100111101, 23'b00000000000000101111101, 23'b00000000000000000000000, 23'b11111111111111111011010, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b00000000000000000001011, 23'b11111111111111100100011, 23'b00000000000001000010011, 23'b11111111111111111110100, 23'b11111111111111111100000, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b11111111111111111110000, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b00000000000000000011010, 23'b11111111111110101110110, 23'b00000000000000001101001, 23'b00000000000000101110111, 23'b11111111111111111111001, 23'b00000000000000011000001, 23'b11111111111111111111111, 23'b00000000000000010011001}, 
{23'b11111111111111001100011, 23'b00000000000000000010010, 23'b11111111111110000100100, 23'b00000000000000000001110, 23'b11111111111111110011001, 23'b11111111111111110101110, 23'b11111111111111111111101, 23'b11111111111111101000101, 23'b11111111111111110110110, 23'b11111111111111101111010, 23'b00000000000000001100000, 23'b00000000000000000110111, 23'b11111111111111010010100, 23'b00000000000000000000001, 23'b11111111111111111111100, 23'b11111111111111111101111, 23'b00000000000000010010000, 23'b11111111111111111010110, 23'b11111111111111111000111, 23'b11111111111111111000100, 23'b11111111111111111111110, 23'b00000000000001000101011, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b11111111111111111101100, 23'b00000000000001010001001, 23'b00000000000000110000010, 23'b00000000000000001000101, 23'b11111111111111100111010, 23'b11111111111111111101011, 23'b00000000000000010000101, 23'b00000000000000001110101}, 
{23'b00000000000000001000101, 23'b00000000000000001010000, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b11111111111110001000000, 23'b00000000000000001011001, 23'b00000000000000000110010, 23'b11111111111111111111111, 23'b00000000000000000000001, 23'b11111111111111010100100, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b11111111111111010110110, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b11111111111110100100111, 23'b00000000000000000010011, 23'b11111111111111111111110, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b00000000000000100001000, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b00000000000001110100101, 23'b00000000000001010111000, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b11111111111111000100001, 23'b00000000000000000000000, 23'b11111111111111111111111}, 
{23'b00000000000000010011011, 23'b00000000000000001101100, 23'b00000000000001000000110, 23'b11111111111111000000011, 23'b00000000000000100001111, 23'b00000000000000011110011, 23'b00000000000000000001100, 23'b00000000000000110001000, 23'b00000000000000000011000, 23'b11111111111111111100111, 23'b00000000000000001001100, 23'b00000000000000000001011, 23'b11111111111111111111110, 23'b00000000000000011110111, 23'b11111111111111111110100, 23'b11111111111111110101110, 23'b00000000000000000000001, 23'b00000000000000001000001, 23'b11111111111111110011101, 23'b00000000000000011001010, 23'b00000000000000001000010, 23'b11111111111101101011011, 23'b11111111111111100010101, 23'b00000000000000010111011, 23'b11111111111111111111111, 23'b11111111111101111110101, 23'b11111111111111011111101, 23'b11111111111111111010000, 23'b11111111111111111111110, 23'b11111111111111110001011, 23'b00000000000000000000000, 23'b11111111111111110101110}, 
{23'b00000000000000000000011, 23'b11111111111111111111111, 23'b11111111111111101000100, 23'b11111111111111010100111, 23'b00000000000000001010101, 23'b00000000000000000000000, 23'b00000000000000011000011, 23'b11111111111111111110100, 23'b00000000000000111111111, 23'b11111111111111111110111, 23'b00000000000000000000000, 23'b11111111111110101000000, 23'b11111111111111111111111, 23'b00000000000000100000001, 23'b11111111111111111111111, 23'b11111111111110111101010, 23'b00000000000000000000000, 23'b11111111111111111101000, 23'b00000000000001000011010, 23'b11111111111111111111111, 23'b11111111111110010000001, 23'b11111111111111111111111, 23'b00000000000001000010000, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b00000000000000100011100, 23'b11111111111111100111111, 23'b00000000000000010001101, 23'b00000000000000000000000, 23'b11111111111111001100011, 23'b00000000000000000000000, 23'b00000000000000000000101}, 
{23'b11111111111111001000101, 23'b00000000000000000000010, 23'b00000000000000000000001, 23'b11111111111111111110011, 23'b00000000000001111110111, 23'b11111111111111100000001, 23'b11111111111111111110100, 23'b11111111111111111110001, 23'b11111111111111110100100, 23'b11111111111111110011000, 23'b00000000000000010000101, 23'b00000000000000100010000, 23'b11111111111111110110100, 23'b00000000000000111111111, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b11111111111110110111010, 23'b11111111111111111111110, 23'b00000000000000000000000, 23'b11111111111111101011100, 23'b00000000000000000000100, 23'b00000000000000001001100, 23'b00000000000000000011011, 23'b11111111111111111101101, 23'b11111111111111110010111, 23'b11111111111111001100000, 23'b11111111111110110100010, 23'b00000000000000000000000, 23'b11111111111111100011000, 23'b00000000000000001010001, 23'b11111111111111111111111, 23'b00000000000000010011010}, 
{23'b11111111111110010110001, 23'b11111111111111010111111, 23'b11111111111111011000000, 23'b00000000000000000000000, 23'b00000000000010010010001, 23'b11111111111111000111000, 23'b00000000000000000000000, 23'b11111111111111110010001, 23'b11111111111110010111000, 23'b00000000000000100011011, 23'b11111111111111111111111, 23'b00000000000010010001001, 23'b00000000000000000000000, 23'b11111111111111110011110, 23'b11111111111111111111111, 23'b00000000000000001000000, 23'b11111111111111111011001, 23'b00000000000000000000000, 23'b11111111111111110100000, 23'b00000000000001111110110, 23'b00000000000000001001111, 23'b11111111111111110101010, 23'b00000000000000011100000, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b11111111111111100111000, 23'b11111111111111110100000, 23'b11111111111110001000001, 23'b11111111111111011011000, 23'b11111111111111111111111, 23'b11111111111111111111101, 23'b11111111111111110000111}, 
{23'b00000000000000111001110, 23'b11111111111100110011010, 23'b11111111111101000110100, 23'b11111111111111010100011, 23'b00000000000010101011010, 23'b11111111111111111111111, 23'b11111111111110100111010, 23'b00000000000001000011110, 23'b00000000000000001111001, 23'b00000000000000000000001, 23'b00000000000000110101010, 23'b11111111111110111010100, 23'b00000000000000000000001, 23'b00000000000000000001000, 23'b11111111111111110111111, 23'b00000000000000000100100, 23'b11111111111111100101011, 23'b11111111111100010100000, 23'b00000000000000101010111, 23'b00000000000001011000010, 23'b00000000000001000011110, 23'b00000000000000000000101, 23'b00000000000000000111011, 23'b11111111111110011000110, 23'b11111111111101011110000, 23'b11111111111111111110101, 23'b11111111111110110011010, 23'b11111111111110001010110, 23'b11111111111111001110000, 23'b11111111111100011111011, 23'b00000000000001101011010, 23'b00000000000001101101111}, 
{23'b00000000000000000000000, 23'b00000000000000000000001, 23'b00000000000000000000100, 23'b00000000000000000000000, 23'b00000000000001000010010, 23'b11111111111111010000001, 23'b00000000000000000100100, 23'b00000000000000010010101, 23'b11111111111110100110101, 23'b00000000000000001001011, 23'b11111111111111111110110, 23'b11111111111111111111110, 23'b11111111111111111111111, 23'b00000000000000111101010, 23'b00000000000000001101010, 23'b00000000000000000101100, 23'b00000000000000001111110, 23'b00000000000001010101010, 23'b11111111111111001000000, 23'b00000000000000000000000, 23'b11111111111111010101111, 23'b11111111111111111111111, 23'b00000000000001010000100, 23'b00000000000000000010000, 23'b11111111111111111111010, 23'b11111111111101110000010, 23'b11111111111111111101101, 23'b11111111111111011000011, 23'b11111111111111110000011, 23'b00000000000000000000111, 23'b00000000000000100010100, 23'b00000000000000011010100}, 
{23'b11111111111111110100111, 23'b00000000000000100010010, 23'b11111111111110110010001, 23'b00000000000000000101010, 23'b00000000000000110001100, 23'b11111111111111110101111, 23'b11111111111111111110110, 23'b00000000000000101001110, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b11111111111111101111010, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b11111111111111110111001, 23'b11111111111111100000110, 23'b11111111111111101111000, 23'b11111111111111110001100, 23'b11111111111111101111111, 23'b11111111111111100011111, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b11111111111111110100100, 23'b11111111111111101110111, 23'b00000000000001100101110, 23'b00000000000000000000000, 23'b11111111111110100011110, 23'b11111111111111111101110, 23'b00000000000000011111100, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b00000000000001000000001, 23'b11111111111111111111111}, 
{23'b11111111111111111111111, 23'b00000000000000000001000, 23'b11111111111111111111111, 23'b11111111111111011000000, 23'b11111111111100100011110, 23'b00000000000000000000001, 23'b00000000000000000000000, 23'b11111111111111111110010, 23'b11111111111101100110100, 23'b00000000000000010100111, 23'b11111111111111100110111, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b11111111111110100001010, 23'b11111111111111110100010, 23'b11111111111111111111111, 23'b00000000000000000000010, 23'b00000000000000000010000, 23'b00000000000000001001010, 23'b00000000000001011000011, 23'b11111111111111100001011, 23'b11111111111110110011011, 23'b00000000000000000000000, 23'b11111111111110111101111, 23'b11111111111111100110101, 23'b11111111111111000100110, 23'b11111111111111111110000, 23'b11111111111111111100110, 23'b11111111111111111011010, 23'b11111111111110000111011, 23'b11111111111111110111010, 23'b00000000000000111110000}, 
{23'b00000000000000011100111, 23'b00000000000000111000000, 23'b11111111111111111111011, 23'b00000000000000101000110, 23'b11111111111111001010000, 23'b11111111111111100000001, 23'b00000000000000011000011, 23'b00000000000000010001100, 23'b11111111111111110011111, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b11111111111110101101111, 23'b11111111111111111111111, 23'b00000000000000100100111, 23'b11111111111111100010101, 23'b00000000000000001000111, 23'b11111111111111111111101, 23'b11111111111111111111101, 23'b00000000000000110101000, 23'b11111111111110101100010, 23'b00000000000001000111111, 23'b00000000000000001100001, 23'b00000000000000000000000, 23'b00000000000000110110001, 23'b00000000000000000000110, 23'b11111111111111110110110, 23'b11111111111110011110100, 23'b11111111111111100011111, 23'b11111111111111010100011, 23'b00000000000000101101011}, 
{23'b00000000000000000000000, 23'b00000000000000000001110, 23'b11111111111110100010010, 23'b11111111111111111111011, 23'b00000000000000110100111, 23'b11111111111111011011110, 23'b11111111111111111100111, 23'b11111111111111111111111, 23'b00000000000000000101001, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b11111111111111001011110, 23'b00000000000000011000100, 23'b00000000000000000001100, 23'b00000000000000000000000, 23'b00000000000000001001100, 23'b11111111111111111111111, 23'b11111111111111011001111, 23'b00000000000000000100100, 23'b00000000000000000000000, 23'b11111111111111110111001, 23'b11111111111111111010011, 23'b00000000000001001011110, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b11111111111110110101000, 23'b11111111111110101100010, 23'b00000000000000111101110, 23'b11111111111111111111101, 23'b11111111111111111111111, 23'b00000000000000000111000, 23'b00000000000001001000010}, 
{23'b11111111111110101000110, 23'b11111111111111111111111, 23'b11111111111111001001100, 23'b00000000000000000001000, 23'b11111111111110100101100, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b11111111111111101111010, 23'b11111111111101110111101, 23'b11111111111111111001011, 23'b00000000000000000000000, 23'b11111111111111111101111, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b11111111111111111101110, 23'b11111111111111110011010, 23'b11111111111111011010001, 23'b11111111111111100111100, 23'b00000000000000010000111, 23'b11111111111111111111011, 23'b11111111111111111001100, 23'b00000000000000000000000, 23'b00000000000001010110001, 23'b11111111111111111111111, 23'b00000000000000100110010, 23'b00000000000000010111011, 23'b11111111111111011100110, 23'b00000000000000110110100, 23'b11111111111111110100010, 23'b00000000000000000000000, 23'b11111111111111111111101, 23'b00000000000010010101000}, 
{23'b11111111111110101111100, 23'b00000000000000000111100, 23'b00000000000000001100111, 23'b11111111111111111000110, 23'b00000000000000111110100, 23'b11111111111110110010101, 23'b11111111111111111110001, 23'b00000000000001000011111, 23'b00000000000000101000110, 23'b00000000000000000010010, 23'b11111111111111111111111, 23'b11111111111111101110011, 23'b11111111111111101001000, 23'b11111111111111101111011, 23'b11111111111111110011010, 23'b00000000000000010111000, 23'b11111111111111111111111, 23'b00000000000000000010000, 23'b00000000000000100100001, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b00000000000000000011110, 23'b00000000000001000000100, 23'b00000000000000001011101, 23'b00000000000000000001101, 23'b11111111111111100100011, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b11111111111111111100011, 23'b11111111111111111100111, 23'b11111111111111111111111, 23'b00000000000000010001010}, 
{23'b11111111111111111111111, 23'b00000000000000000000111, 23'b11111111111111001001101, 23'b11111111111111101100111, 23'b00000000000001001000001, 23'b11111111111111111111111, 23'b11111111111111101100001, 23'b00000000000000111110100, 23'b11111111111111110010011, 23'b00000000000001001010101, 23'b00000000000000010101111, 23'b11111111111111100001001, 23'b00000000000000000000001, 23'b00000000000000000000111, 23'b11111111111111111100001, 23'b00000000000000000101011, 23'b11111111111111101100010, 23'b11111111111110111100100, 23'b00000000000001000111001, 23'b00000000000000100111110, 23'b00000000000010100010011, 23'b00000000000000110011011, 23'b00000000000000111111100, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b00000000000000001110101, 23'b00000000000000010100010, 23'b11111111111110010100011, 23'b11111111111111111111111, 23'b11111111111111111110101, 23'b11111111111111111110010}, 
{23'b00000000000000000000001, 23'b11111111111111101001100, 23'b11111111111111100101011, 23'b00000000000000000000000, 23'b11111111111111000001101, 23'b00000000000000000000000, 23'b00000000000000110001000, 23'b00000000000000011011111, 23'b00000000000000001101100, 23'b11111111111111100110101, 23'b00000000000000000000000, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b11111111111111110101000, 23'b00000000000000110011101, 23'b11111111111111111111111, 23'b11111111111111111111110, 23'b11111111111110110010100, 23'b00000000000000000000000, 23'b11111111111111001110101, 23'b11111111111111111111101, 23'b00000000000000000000000, 23'b11111111111111111110111, 23'b00000000000000000011110, 23'b00000000000000000100011, 23'b00000000000000000111001, 23'b00000000000000100011011, 23'b11111111111111101111010, 23'b11111111111111111110000, 23'b11111111111110001101001, 23'b00000000000000010100001}, 
{23'b00000000000001110001000, 23'b11111111111111111101110, 23'b00000000000000010000111, 23'b11111111111111100101001, 23'b11111111111111101010001, 23'b00000000000000001000100, 23'b00000000000000101001000, 23'b00000000000000000000000, 23'b00000000000010000110111, 23'b00000000000000000000000, 23'b11111111111111111010100, 23'b00000000000000000100110, 23'b00000000000000011000000, 23'b11111111111111111111010, 23'b00000000000000001101101, 23'b00000000000000011010011, 23'b11111111111111111110111, 23'b11111111111110001110000, 23'b11111111111111110001100, 23'b11111111111111111111100, 23'b00000000000000011101110, 23'b00000000000000000000011, 23'b11111111111111111111111, 23'b00000000000000011100110, 23'b00000000000000000100100, 23'b11111111111110111100100, 23'b11111111111111100101101, 23'b00000000000000100001110, 23'b11111111111111111000110, 23'b00000000000001000010000, 23'b11111111111111111111101, 23'b11111111111111010010001}, 
{23'b00000000000000000011010, 23'b00000000000000011010000, 23'b11111111111111111111111, 23'b11111111111111110110000, 23'b11111111111110100101101, 23'b11111111111111111111111, 23'b00000000000000001011110, 23'b11111111111111110100001, 23'b00000000000000101010001, 23'b11111111111111110111010, 23'b11111111111111111111110, 23'b11111111111111110111011, 23'b11111111111111111111111, 23'b11111111111111110110100, 23'b00000000000000000000000, 23'b00000000000001010000001, 23'b00000000000000000000000, 23'b11111111111111111111100, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b00000000000000001000101, 23'b00000000000000100000001, 23'b00000000000000000000000, 23'b00000000000000000001000, 23'b00000000000000001000010, 23'b11111111111111111111110, 23'b00000000000000000000000, 23'b00000000000000000101001, 23'b00000000000000000000011, 23'b00000000000000011000110}, 
{23'b11111111111110110000111, 23'b00000000000000100001010, 23'b00000000000000000100100, 23'b11111111111111100101000, 23'b11111111111110011001110, 23'b11111111111111111011010, 23'b00000000000000010001001, 23'b11111111111110011010010, 23'b00000000000010000010111, 23'b00000000000000010010010, 23'b00000000000000000100000, 23'b00000000000000011000001, 23'b00000000000000001011010, 23'b00000000000000000000001, 23'b00000000000001101000011, 23'b11111111111111101010011, 23'b00000000000000000001010, 23'b00000000000000000000000, 23'b11111111111111111110010, 23'b00000000000000000000111, 23'b11111111111110010001011, 23'b00000000000000000100010, 23'b00000000000000100111001, 23'b00000000000000001001100, 23'b00000000000000001001001, 23'b11111111111101010111111, 23'b11111111111110101000101, 23'b11111111111111000010011, 23'b00000000000000000000101, 23'b11111111111111111111100, 23'b00000000000001010011011, 23'b11111111111111001011100}, 
{23'b11111111111111111100101, 23'b11111111111111001110001, 23'b11111111111111100101100, 23'b11111111111110010111011, 23'b11111111111110111101011, 23'b00000000000001010110000, 23'b00000000000001001111010, 23'b11111111111111010100011, 23'b00000000000000001010101, 23'b11111111111111110110000, 23'b11111111111111100111111, 23'b11111111111110111111101, 23'b00000000000000011010011, 23'b11111111111110110111010, 23'b00000000000000110000010, 23'b11111111111111111111111, 23'b00000000000001010101111, 23'b11111111111111111111111, 23'b11111111111111111110000, 23'b11111111111111011101010, 23'b11111111111111110101010, 23'b11111111111111101111011, 23'b11111111111110111011111, 23'b00000000000000010101000, 23'b11111111111111111111111, 23'b11111111111111111110011, 23'b11111111111111000101100, 23'b00000000000001010000100, 23'b00000000000001000111011, 23'b11111111111111101000110, 23'b11111111111101011110100, 23'b00000000000000100100100}, 
{23'b00000000000000000000000, 23'b11111111111111111001011, 23'b11111111111111111111111, 23'b11111111111111100111000, 23'b00000000000000000111010, 23'b00000000000000000010010, 23'b00000000000000010001110, 23'b00000000000000000001011, 23'b00000000000000011110001, 23'b11111111111111111111110, 23'b00000000000000000000000, 23'b00000000000000011000011, 23'b00000000000000000000011, 23'b00000000000000000011001, 23'b11111111111111011110000, 23'b11111111111111100100011, 23'b00000000000000000000000, 23'b00000000000000101110100, 23'b00000000000000001110100, 23'b00000000000000100000001, 23'b11111111111111111011110, 23'b11111111111111010111000, 23'b11111111111111111111111, 23'b00000000000000010011000, 23'b11111111111111111111111, 23'b00000000000000001000010, 23'b11111111111111111110110, 23'b00000000000000010001010, 23'b00000000000000000000000, 23'b00000000000000010101010, 23'b11111111111110011110110, 23'b11111111111111111111111}, 
{23'b00000000000001001111011, 23'b11111111111111111101101, 23'b00000000000000100110011, 23'b11111111111110110001110, 23'b11111111111111001110100, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b00000000000000000111000, 23'b00000000000000000000100, 23'b11111111111111011111110, 23'b00000000000000000000000, 23'b00000000000000000000100, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b11111111111111011110111, 23'b00000000000000100100100, 23'b11111111111111111111100, 23'b11111111111111111000000, 23'b00000000000000000000000, 23'b00000000000000011110101, 23'b11111111111111001100100, 23'b00000000000000011101101, 23'b00000000000000100011110, 23'b00000000000000100001000, 23'b11111111111111111111111, 23'b00000000000010001101001, 23'b11111111111111011000110, 23'b00000000000001011101000, 23'b11111111111111110010110, 23'b11111111111110100011101, 23'b11111111111111010011100, 23'b00000000000000100011101}, 
{23'b11111111111101110100111, 23'b11111111111111111001001, 23'b11111111111111011000100, 23'b11111111111111111111111, 23'b00000000000001000010110, 23'b11111111111111010010010, 23'b11111111111111110000101, 23'b00000000000000111100111, 23'b00000000000000011000001, 23'b11111111111111000011000, 23'b00000000000000000000000, 23'b11111111111111111000110, 23'b11111111111111111101011, 23'b00000000000000100011001, 23'b11111111111111000001000, 23'b11111111111111111101001, 23'b00000000000000000000000, 23'b11111111111111111111110, 23'b11111111111111111011111, 23'b00000000000000000000000, 23'b11111111111111001111010, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b11111111111110101011111, 23'b00000000000000010001111, 23'b00000000000010011110101, 23'b00000000000001011000100, 23'b11111111111111110110110, 23'b11111111111111010110111, 23'b11111111111110001101001, 23'b00000000000000000000000, 23'b11111111111111110011100}, 
{23'b00000000000000000101011, 23'b00000000000000110110101, 23'b00000000000000000101011, 23'b11111111111111011001010, 23'b00000000000000000001001, 23'b11111111111111111001011, 23'b00000000000000000000000, 23'b00000000000000110101010, 23'b00000000000000110111000, 23'b11111111111111011101110, 23'b00000000000000100011111, 23'b00000000000000000110001, 23'b11111111111111111111111, 23'b11111111111111111100010, 23'b11111111111111010111010, 23'b00000000000001000000110, 23'b11111111111111110101001, 23'b11111111111110101101010, 23'b00000000000000011101010, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b00000000000000011101111, 23'b11111111111111101100111, 23'b11111111111111111110110, 23'b11111111111111110010110, 23'b00000000000000010110100, 23'b11111111111111011100000, 23'b00000000000000100010010, 23'b11111111111110100010111, 23'b00000000000000010100100, 23'b11111111111111111111111, 23'b00000000000000101000000}, 
{23'b11111111111111110101000, 23'b00000000000000000000001, 23'b00000000000000010110110, 23'b00000000000000000000000, 23'b11111111111111110000011, 23'b11111111111111111111010, 23'b00000000000000011010010, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b00000000000000000001010, 23'b00000000000000000000000, 23'b00000000000000000101000, 23'b11111111111111100100110, 23'b00000000000000000010101, 23'b00000000000000011100010, 23'b00000000000000001011111, 23'b00000000000000011011000, 23'b11111111111111111111110, 23'b11111111111111111111101, 23'b00000000000000100000110, 23'b00000000000000111111010, 23'b11111111111111100110111, 23'b00000000000000000000000, 23'b11111111111111111111011, 23'b00000000000000000010111, 23'b11111111111110001001111, 23'b11111111111111111111110, 23'b11111111111111101101111, 23'b11111111111111111111111, 23'b00000000000010010000100, 23'b00000000000000000000000, 23'b11111111111111001011010}, 
{23'b11111111111111111001001, 23'b11111111111111100001011, 23'b11111111111111111101101, 23'b00000000000000000001110, 23'b00000000000000010111001, 23'b11111111111111111111111, 23'b00000000000000000000000, 23'b11111111111111111010000, 23'b00000000000000010010000, 23'b11111111111111111101111, 23'b00000000000000000000000, 23'b00000000000000001000000, 23'b00000000000001001011100, 23'b11111111111111100101111, 23'b00000000000000000011001, 23'b11111111111100100110110, 23'b11111111111111111101001, 23'b11111111111111110000100, 23'b00000000000000000010000, 23'b11111111111111110011001, 23'b00000000000000010111100, 23'b11111111111111000110101, 23'b00000000000000011101001, 23'b00000000000000011010111, 23'b11111111111111111100101, 23'b11111111111101001001111, 23'b11111111111111000101011, 23'b11111111111111111010011, 23'b11111111111111111011010, 23'b00000000000001100011111, 23'b11111111111111111110100, 23'b00000000000000100111011}, 
{23'b00000000000000001100000, 23'b00000000000000000000000, 23'b00000000000000101100100, 23'b11111111111111100010111, 23'b11111111111111101110011, 23'b00000000000000111100111, 23'b11111111111111010111000, 23'b00000000000000001110101, 23'b11111111111110110000110, 23'b00000000000000000010001, 23'b00000000000000000100010, 23'b11111111111111101010100, 23'b00000000000000000000001, 23'b00000000000000000000000, 23'b11111111111111001111111, 23'b00000000000001101110101, 23'b11111111111111000000110, 23'b11111111111111111100111, 23'b00000000000000011110011, 23'b11111111111111111111111, 23'b00000000000000010001101, 23'b11111111111110000101010, 23'b00000000000001010000001, 23'b11111111111111111111111, 23'b11111111111111100000010, 23'b00000000000001111100000, 23'b00000000000000100101011, 23'b11111111111111010111100, 23'b11111111111111011101100, 23'b11111111111101110110011, 23'b11111111111111111101011, 23'b00000000000000000100000}, 
{23'b11111111111111111111111, 23'b00000000000000000001101, 23'b11111111111111110111000, 23'b11111111111110111011011, 23'b11111111111111111111111, 23'b11111111111110011011100, 23'b00000000000000000000000, 23'b00000000000001001101101, 23'b00000000000000111110100, 23'b00000000000000000100110, 23'b00000000000000000000000, 23'b11111111111111100011110, 23'b00000000000001010101000, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b00000000000001101111000, 23'b00000000000000000000011, 23'b11111111111111110101110, 23'b11111111111111110010111, 23'b11111111111110101101100, 23'b00000000000000100001101, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b00000000000000001000000, 23'b11111111111111101101110, 23'b11111111111110001010000, 23'b00000000000001000110101, 23'b11111111111110001110011, 23'b00000000000000001101000, 23'b11111111111111101011110, 23'b00000000000000000000000}, 
{23'b00000000000000001111101, 23'b00000000000000101111101, 23'b00000000000000000010011, 23'b11111111111111111111001, 23'b11111111111110001010011, 23'b00000000000000000000001, 23'b11111111111111111111111, 23'b00000000000000111110000, 23'b00000000000001000110111, 23'b11111111111111111111111, 23'b11111111111111111111111, 23'b11111111111111111111101, 23'b00000000000000000000000, 23'b00000000000000000000100, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b00000000000000000000000, 23'b11111111111111111111110, 23'b00000000000000101011100, 23'b11111111111111100101101, 23'b11111111111110010001011, 23'b11111111111111110111100, 23'b11111111111111100110101, 23'b11111111111111100111111, 23'b11111111111111101110010, 23'b11111111111111111111110, 23'b11111111111111101111111, 23'b11111111111111111010011, 23'b11111111111111111101010, 23'b00000000000000100100001, 23'b11111111111111111111111, 23'b00000000000001110110101}
};

localparam logic signed [22:0] bias [32] = '{
23'b00000000000101111001011,  // 1.474280834197998
23'b00000000000010110001000,  // 0.6914801001548767
23'b00000000000101110000110,  // 1.4406442642211914
23'b00000000000101101000011,  // 1.408045768737793
23'b00000000000011111100100,  // 0.9864811301231384
23'b00000000000011011101000,  // 0.8636202812194824
23'b11111111111101100010011,  // -0.6153604388237
23'b00000000000001111011111,  // 0.4839226007461548
23'b00000000000001111100011,  // 0.4862793982028961
23'b00000000000001011111001,  // 0.37162142992019653
23'b00000000000001110101101,  // 0.45989668369293213
23'b00000000000101001100110,  // 1.2998151779174805
23'b11111111111011111011110,  // -1.016528844833374
23'b11111111111110100101110,  // -0.35249894857406616
23'b00000000000001110010001,  // 0.44582197070121765
23'b11111111111111100011010,  // -0.1119980737566948
23'b11111111111111101110110,  // -0.06717441976070404
23'b00000000000000000001001,  // 0.00487547367811203
23'b00000000000000110001110,  // 0.1946917623281479
23'b11111111111100111000011,  // -0.7796769738197327
23'b00000000000010111010100,  // 0.7287401556968689
23'b00000000000110110111000,  // 1.714877724647522
23'b11111111111001100111001,  // -1.5971007347106934
23'b00000000000000010010111,  // 0.07393483817577362
23'b00000000000001010010100,  // 0.3225609362125397
23'b00000000000011011000011,  // 0.8453295230865479
23'b00000000000011100110000,  // 0.898597240447998
23'b00000000000001000001001,  // 0.2548799514770508
23'b00000000000011111001001,  // 0.9735668301582336
23'b00000000000100100000010,  // 1.1261906623840332
23'b00000000000001110010100,  // 0.44768181443214417
23'b11111111110110100001111   // -2.3676068782806396
};
endpackage