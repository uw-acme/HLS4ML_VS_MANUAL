// Width: 22
// NFRAC: 11
package dense_4_22_11;

localparam logic signed [21:0] weights [32][5] = '{ 
{22'b1111111111111111100111, 22'b0000000000001010000110, 22'b1111111111110110011101, 22'b0000000000000010000110, 22'b1111111111111100100110}, 
{22'b1111111111101110001001, 22'b1111111111111110001111, 22'b0000000000001110101110, 22'b1111111111111111100110, 22'b0000000000000000100010}, 
{22'b0000000000001011111000, 22'b0000000000000110110001, 22'b1111111111111111000110, 22'b1111111111110011000001, 22'b1111111111111001010000}, 
{22'b1111111111110011111110, 22'b1111111111110100000100, 22'b1111111111111100011011, 22'b0000000000001001110110, 22'b0000000000000111100001}, 
{22'b0000000000000011111010, 22'b0000000000000100000111, 22'b0000000000000101000001, 22'b1111111111111111011010, 22'b1111111111011111100101}, 
{22'b0000000000001010011101, 22'b1111111111110011011000, 22'b0000000000000101110011, 22'b1111111111111010110101, 22'b1111111111111010100011}, 
{22'b1111111111110011001010, 22'b0000000000000001001000, 22'b1111111111111111111111, 22'b0000000000000101100100, 22'b0000000000000010001101}, 
{22'b1111111111111111111100, 22'b0000000000001001000110, 22'b1111111111110011011101, 22'b0000000000000101001101, 22'b0000000000000100010110}, 
{22'b0000000000000101001110, 22'b1111111111111010100101, 22'b0000000000000000000010, 22'b1111111111110001001110, 22'b1111111111111000000010}, 
{22'b1111111111111111111111, 22'b1111111111110111011110, 22'b0000000000000101101100, 22'b0000000000001101110000, 22'b0000000000000000000000}, 
{22'b1111111111111011110101, 22'b1111111111111011010111, 22'b0000000000000000000000, 22'b0000000000010010100110, 22'b1111111111110111011011}, 
{22'b0000000000000101011010, 22'b0000000000000111010101, 22'b1111111111110101000111, 22'b1111111111111111000111, 22'b0000000000000011111001}, 
{22'b0000000000000000000000, 22'b0000000000000101010111, 22'b0000000000000000010010, 22'b1111111111111001010110, 22'b1111111111101100000100}, 
{22'b0000000000000101101011, 22'b0000000000000010000010, 22'b0000000000001101011011, 22'b1111111111111101110000, 22'b1111111111110010010011}, 
{22'b0000000000000010111001, 22'b1111111111111110011101, 22'b1111111111110100011101, 22'b1111111111111110111100, 22'b0000000000010001001010}, 
{22'b1111111111110000110101, 22'b1111111111111000001011, 22'b1111111111111000111000, 22'b0000000000001100110000, 22'b0000000000000001000001}, 
{22'b0000000000001011000100, 22'b1111111111111010100000, 22'b1111111111111011101010, 22'b1111111111111000110001, 22'b1111111111111110000101}, 
{22'b0000000000000110001111, 22'b1111111111111110101101, 22'b1111111111110010110011, 22'b1111111111111111000001, 22'b0000000000000010010000}, 
{22'b0000000000001000010001, 22'b0000000000000001010101, 22'b1111111111111001000001, 22'b0000000000000000000000, 22'b1111111111110011111110}, 
{22'b0000000000000111011001, 22'b1111111111111101001110, 22'b1111111111111001001100, 22'b0000000000000110101000, 22'b0000000000000011000010}, 
{22'b0000000000000010001010, 22'b1111111111111111000001, 22'b0000000000001001100001, 22'b1111111111110010001101, 22'b1111111111111111010100}, 
{22'b0000000000000000000000, 22'b0000000000000011110001, 22'b0000000000001111100100, 22'b1111111111101111011010, 22'b1111111111101100001111}, 
{22'b1111111111111100110110, 22'b0000000000000011100000, 22'b0000000000000101101010, 22'b1111111111110100100101, 22'b0000000000010000101101}, 
{22'b1111111111111111111111, 22'b0000000000000101010001, 22'b0000000000001001000010, 22'b0000000000000001001101, 22'b1111111111101101101100}, 
{22'b1111111111111010100101, 22'b0000000000001011101010, 22'b1111111111111000110110, 22'b0000000000000000001011, 22'b0000000000001100011010}, 
{22'b0000000000000000110101, 22'b0000000000001000100000, 22'b0000000000000000111100, 22'b1111111111101000000100, 22'b0000000000010001100010}, 
{22'b1111111111110001010010, 22'b1111111111111000001101, 22'b0000000000000110110110, 22'b0000000000000111110100, 22'b0000000000000110011101}, 
{22'b0000000000000000001000, 22'b0000000000000111101101, 22'b1111111111111110110101, 22'b1111111111111011001011, 22'b0000000000000001000000}, 
{22'b1111111111111100101010, 22'b0000000000000111111000, 22'b1111111111101111111000, 22'b0000000000000100011100, 22'b1111111111111010111011}, 
{22'b1111111111111111011010, 22'b0000000000000100100001, 22'b1111111111111010100110, 22'b1111111111110011001011, 22'b0000000000010010111111}, 
{22'b0000000000001110010111, 22'b0000000000000010001111, 22'b0000000000001010011000, 22'b1111111111101101001000, 22'b1111111111110101111010}, 
{22'b1111111111111110000110, 22'b1111111111110011101001, 22'b0000000000001011101101, 22'b0000000000000010010001, 22'b0000000000000100000101}
};

localparam logic signed [21:0] bias [5] = '{
22'b1111111111111110000000,  // -0.06223141402006149
22'b1111111111111101111111,  // -0.06270556896924973
22'b1111111111111101110000,  // -0.07014333456754684
22'b0000000000000010101000,  // 0.0820775106549263
22'b0000000000000110111001   // 0.2155742198228836
};
endpackage