// Width: 6
// NFRAC: 3
package dense_1_6_3;

localparam logic signed [5:0] weights [16][64] = '{ 
{6'b000010, 6'b111010, 6'b111110, 6'b111110, 6'b111100, 6'b000000, 6'b110111, 6'b000000, 6'b000000, 6'b000010, 6'b000000, 6'b111100, 6'b111111, 6'b000001, 6'b000000, 6'b111101, 6'b000001, 6'b000000, 6'b000000, 6'b111111, 6'b000011, 6'b111101, 6'b111111, 6'b000011, 6'b111101, 6'b111010, 6'b111101, 6'b111110, 6'b111111, 6'b111111, 6'b000000, 6'b000001, 6'b000001, 6'b111111, 6'b000000, 6'b000010, 6'b111111, 6'b111101, 6'b000000, 6'b000001, 6'b111111, 6'b000010, 6'b111101, 6'b000111, 6'b111111, 6'b000011, 6'b000000, 6'b000001, 6'b000001, 6'b111111, 6'b000000, 6'b000001, 6'b000001, 6'b000000, 6'b111111, 6'b111101, 6'b000100, 6'b111100, 6'b000011, 6'b111101, 6'b000110, 6'b111111, 6'b000000, 6'b000000}, 
{6'b000000, 6'b111101, 6'b111110, 6'b111101, 6'b111101, 6'b000000, 6'b111001, 6'b111111, 6'b111110, 6'b000001, 6'b000000, 6'b111111, 6'b000001, 6'b000000, 6'b111111, 6'b000001, 6'b111111, 6'b000000, 6'b111110, 6'b111101, 6'b000011, 6'b111111, 6'b000000, 6'b000101, 6'b000010, 6'b111110, 6'b111110, 6'b111111, 6'b111111, 6'b111100, 6'b111111, 6'b000011, 6'b000010, 6'b000100, 6'b000101, 6'b000000, 6'b111111, 6'b111100, 6'b000000, 6'b000001, 6'b000000, 6'b000001, 6'b111110, 6'b000010, 6'b000001, 6'b000000, 6'b111101, 6'b000000, 6'b000010, 6'b000000, 6'b000000, 6'b001001, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b000010, 6'b111101, 6'b000111, 6'b000000, 6'b000100, 6'b000001, 6'b000110, 6'b000001}, 
{6'b111111, 6'b000000, 6'b111111, 6'b111110, 6'b111110, 6'b000000, 6'b001011, 6'b111111, 6'b110101, 6'b111111, 6'b111111, 6'b111111, 6'b111110, 6'b000000, 6'b111111, 6'b000001, 6'b000111, 6'b111111, 6'b000000, 6'b000000, 6'b000011, 6'b111010, 6'b000100, 6'b111010, 6'b000111, 6'b111101, 6'b111110, 6'b111010, 6'b001010, 6'b000010, 6'b000000, 6'b000100, 6'b001000, 6'b110110, 6'b111111, 6'b000000, 6'b111110, 6'b000111, 6'b111111, 6'b000010, 6'b000010, 6'b000010, 6'b111111, 6'b111111, 6'b111111, 6'b000001, 6'b111101, 6'b111110, 6'b111111, 6'b000011, 6'b111110, 6'b000001, 6'b111111, 6'b000001, 6'b111110, 6'b111111, 6'b111101, 6'b111010, 6'b111111, 6'b000000, 6'b001100, 6'b000000, 6'b111111, 6'b111101}, 
{6'b111100, 6'b111101, 6'b111010, 6'b000010, 6'b111101, 6'b110101, 6'b111111, 6'b111101, 6'b000001, 6'b111111, 6'b001010, 6'b111111, 6'b111001, 6'b000100, 6'b000000, 6'b111111, 6'b111100, 6'b111111, 6'b000000, 6'b111110, 6'b110110, 6'b111111, 6'b111010, 6'b000001, 6'b111100, 6'b111000, 6'b000010, 6'b000101, 6'b001010, 6'b111100, 6'b111011, 6'b000000, 6'b000100, 6'b111001, 6'b111101, 6'b000000, 6'b111010, 6'b000001, 6'b111100, 6'b000000, 6'b000011, 6'b000001, 6'b000000, 6'b000000, 6'b000100, 6'b111110, 6'b111111, 6'b111101, 6'b111111, 6'b111111, 6'b111011, 6'b000000, 6'b111111, 6'b000001, 6'b000010, 6'b000101, 6'b111000, 6'b111000, 6'b111010, 6'b000110, 6'b001101, 6'b111000, 6'b111111, 6'b000011}, 
{6'b000010, 6'b111011, 6'b111101, 6'b111111, 6'b111110, 6'b000010, 6'b000001, 6'b111111, 6'b111011, 6'b111110, 6'b111101, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b000010, 6'b000001, 6'b111100, 6'b000000, 6'b000000, 6'b000001, 6'b111111, 6'b000000, 6'b111111, 6'b001000, 6'b111110, 6'b111101, 6'b111100, 6'b000000, 6'b000001, 6'b000000, 6'b000010, 6'b111111, 6'b000000, 6'b000001, 6'b111111, 6'b000000, 6'b000111, 6'b111101, 6'b111111, 6'b000011, 6'b000001, 6'b111100, 6'b000000, 6'b110111, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b000001, 6'b111111, 6'b000010, 6'b111110, 6'b111010, 6'b111100, 6'b111011, 6'b111011, 6'b000101, 6'b001010, 6'b000110, 6'b000000, 6'b111111}, 
{6'b111100, 6'b111010, 6'b000000, 6'b000010, 6'b000010, 6'b111110, 6'b000100, 6'b111111, 6'b000001, 6'b111111, 6'b111111, 6'b111111, 6'b111110, 6'b000100, 6'b111111, 6'b000000, 6'b111011, 6'b111101, 6'b000000, 6'b111111, 6'b111111, 6'b111101, 6'b111101, 6'b000011, 6'b111101, 6'b111111, 6'b000010, 6'b111111, 6'b111000, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b000001, 6'b000010, 6'b000000, 6'b111111, 6'b111101, 6'b111111, 6'b111110, 6'b111011, 6'b000011, 6'b000000, 6'b000100, 6'b000000, 6'b111111, 6'b000000, 6'b111100, 6'b000001, 6'b000000, 6'b111111, 6'b111101, 6'b000011, 6'b111111, 6'b000010, 6'b000001, 6'b000001, 6'b111111, 6'b111111, 6'b111001, 6'b111110, 6'b111111, 6'b111111}, 
{6'b111101, 6'b111101, 6'b111100, 6'b111111, 6'b111110, 6'b000000, 6'b111010, 6'b111110, 6'b111110, 6'b111111, 6'b111101, 6'b000010, 6'b000000, 6'b000001, 6'b000010, 6'b000000, 6'b000110, 6'b000000, 6'b000001, 6'b000010, 6'b111110, 6'b000010, 6'b111110, 6'b111011, 6'b000001, 6'b000100, 6'b111111, 6'b000000, 6'b111000, 6'b000010, 6'b000010, 6'b111101, 6'b000011, 6'b000101, 6'b000000, 6'b000010, 6'b111111, 6'b000010, 6'b000001, 6'b000000, 6'b111111, 6'b111101, 6'b000001, 6'b000011, 6'b000100, 6'b111110, 6'b111111, 6'b111110, 6'b111110, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000001, 6'b111110, 6'b000110, 6'b000010, 6'b111111, 6'b000011, 6'b000001, 6'b110010, 6'b111011, 6'b111110, 6'b111111}, 
{6'b000000, 6'b000001, 6'b111111, 6'b111111, 6'b111101, 6'b111111, 6'b111101, 6'b000000, 6'b000000, 6'b000011, 6'b000000, 6'b111100, 6'b111111, 6'b000000, 6'b111111, 6'b111100, 6'b111001, 6'b111111, 6'b111011, 6'b111100, 6'b111100, 6'b000010, 6'b000000, 6'b111110, 6'b111100, 6'b000001, 6'b000000, 6'b000011, 6'b000110, 6'b111111, 6'b000000, 6'b000001, 6'b111010, 6'b111101, 6'b000000, 6'b000000, 6'b111101, 6'b000001, 6'b000001, 6'b111110, 6'b111100, 6'b111111, 6'b000000, 6'b111110, 6'b000000, 6'b000001, 6'b111111, 6'b000000, 6'b000000, 6'b111110, 6'b111100, 6'b000011, 6'b000001, 6'b111110, 6'b000001, 6'b111111, 6'b111100, 6'b111110, 6'b111111, 6'b111111, 6'b000110, 6'b000001, 6'b111111, 6'b111111}, 
{6'b000000, 6'b000100, 6'b111011, 6'b111110, 6'b000010, 6'b111110, 6'b001001, 6'b111101, 6'b111111, 6'b000010, 6'b000010, 6'b111111, 6'b111111, 6'b111100, 6'b000010, 6'b000001, 6'b111110, 6'b111111, 6'b000000, 6'b000000, 6'b000010, 6'b111100, 6'b000011, 6'b000100, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b000101, 6'b000000, 6'b111101, 6'b000000, 6'b000011, 6'b111001, 6'b111011, 6'b000001, 6'b000001, 6'b111011, 6'b111110, 6'b111110, 6'b000011, 6'b000011, 6'b000000, 6'b111101, 6'b000000, 6'b000011, 6'b111111, 6'b111111, 6'b000000, 6'b000001, 6'b111111, 6'b111110, 6'b000010, 6'b111110, 6'b000010, 6'b000100, 6'b000000, 6'b000010, 6'b111100, 6'b111101, 6'b000110, 6'b111110, 6'b000000, 6'b111111}, 
{6'b000000, 6'b111100, 6'b000010, 6'b111101, 6'b111111, 6'b000001, 6'b111011, 6'b000001, 6'b000011, 6'b000001, 6'b000010, 6'b000010, 6'b111101, 6'b111111, 6'b111111, 6'b000000, 6'b111000, 6'b000010, 6'b111111, 6'b000000, 6'b111101, 6'b000000, 6'b000001, 6'b111111, 6'b111100, 6'b111111, 6'b111111, 6'b001001, 6'b111010, 6'b000000, 6'b000000, 6'b111111, 6'b111110, 6'b000000, 6'b111111, 6'b111110, 6'b111110, 6'b111110, 6'b111111, 6'b111101, 6'b000010, 6'b000000, 6'b000011, 6'b000000, 6'b000000, 6'b111101, 6'b000000, 6'b111111, 6'b111111, 6'b000001, 6'b000001, 6'b000010, 6'b111111, 6'b111101, 6'b000000, 6'b000000, 6'b000010, 6'b111110, 6'b111011, 6'b000100, 6'b111101, 6'b001001, 6'b111111, 6'b111101}, 
{6'b111011, 6'b111111, 6'b111100, 6'b000001, 6'b000010, 6'b111111, 6'b000100, 6'b111110, 6'b111100, 6'b111101, 6'b111101, 6'b111100, 6'b111110, 6'b000001, 6'b000000, 6'b000000, 6'b000110, 6'b111111, 6'b111111, 6'b000011, 6'b000010, 6'b111011, 6'b111100, 6'b000001, 6'b111100, 6'b111111, 6'b111101, 6'b111101, 6'b111100, 6'b000010, 6'b000001, 6'b111110, 6'b111111, 6'b111000, 6'b111110, 6'b000000, 6'b111110, 6'b111101, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b111010, 6'b000000, 6'b000000, 6'b000010, 6'b111111, 6'b000011, 6'b111110, 6'b000010, 6'b111111, 6'b000001, 6'b111100, 6'b111111, 6'b000100, 6'b000010, 6'b000010, 6'b000000, 6'b111100, 6'b111101, 6'b111010, 6'b111111, 6'b000000}, 
{6'b000010, 6'b000000, 6'b000001, 6'b111111, 6'b000001, 6'b111110, 6'b000001, 6'b000000, 6'b000001, 6'b000010, 6'b111101, 6'b111111, 6'b111111, 6'b111111, 6'b111010, 6'b111101, 6'b000101, 6'b111111, 6'b111111, 6'b000000, 6'b111100, 6'b000000, 6'b000010, 6'b000000, 6'b000000, 6'b000010, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b111110, 6'b111010, 6'b000010, 6'b000010, 6'b111111, 6'b111110, 6'b000000, 6'b111010, 6'b111111, 6'b111111, 6'b000001, 6'b111110, 6'b111111, 6'b000110, 6'b000011, 6'b111111, 6'b111111, 6'b111111, 6'b111110, 6'b000001, 6'b000001, 6'b000001, 6'b000001, 6'b000011, 6'b000010, 6'b000101, 6'b111110, 6'b000011, 6'b000001, 6'b111101, 6'b000000, 6'b111100, 6'b111100, 6'b111100}, 
{6'b000000, 6'b000001, 6'b111110, 6'b000000, 6'b111111, 6'b111111, 6'b111010, 6'b111111, 6'b000010, 6'b000001, 6'b000001, 6'b111100, 6'b111111, 6'b000010, 6'b111111, 6'b000000, 6'b111001, 6'b111111, 6'b000010, 6'b000000, 6'b000001, 6'b111111, 6'b000001, 6'b000011, 6'b111101, 6'b111101, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b000010, 6'b111010, 6'b000010, 6'b000100, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b111101, 6'b111111, 6'b000001, 6'b000101, 6'b111001, 6'b111100, 6'b000001, 6'b111111, 6'b000011, 6'b111110, 6'b111101, 6'b111101, 6'b111111, 6'b000000, 6'b111110, 6'b111001, 6'b111110, 6'b111111, 6'b000000, 6'b111011, 6'b001000, 6'b111011, 6'b000100, 6'b000001}, 
{6'b000000, 6'b111110, 6'b000101, 6'b111101, 6'b111100, 6'b000000, 6'b000010, 6'b000010, 6'b111110, 6'b111110, 6'b000000, 6'b000001, 6'b000001, 6'b000000, 6'b111110, 6'b000001, 6'b000011, 6'b111111, 6'b111101, 6'b000000, 6'b000000, 6'b000000, 6'b111101, 6'b000000, 6'b000110, 6'b000000, 6'b000001, 6'b111001, 6'b111111, 6'b000000, 6'b111110, 6'b111101, 6'b000011, 6'b111111, 6'b111111, 6'b111101, 6'b000001, 6'b000010, 6'b111111, 6'b111111, 6'b111110, 6'b000001, 6'b000000, 6'b111010, 6'b000010, 6'b000011, 6'b111111, 6'b000000, 6'b111100, 6'b111111, 6'b111111, 6'b111101, 6'b000000, 6'b111110, 6'b000000, 6'b111001, 6'b111111, 6'b111111, 6'b000010, 6'b000100, 6'b111010, 6'b000100, 6'b000000, 6'b111111}, 
{6'b000010, 6'b001001, 6'b000011, 6'b000010, 6'b111100, 6'b111101, 6'b101011, 6'b111100, 6'b000011, 6'b111111, 6'b000010, 6'b000110, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b111110, 6'b111110, 6'b000001, 6'b111011, 6'b111010, 6'b111111, 6'b111011, 6'b000000, 6'b101101, 6'b000110, 6'b000111, 6'b000100, 6'b110010, 6'b111101, 6'b111010, 6'b111001, 6'b101011, 6'b000101, 6'b111111, 6'b000010, 6'b000000, 6'b110100, 6'b000000, 6'b000000, 6'b000000, 6'b001000, 6'b111110, 6'b111010, 6'b000111, 6'b111100, 6'b111101, 6'b111100, 6'b000011, 6'b000100, 6'b111111, 6'b111101, 6'b111111, 6'b111111, 6'b000000, 6'b111100, 6'b000100, 6'b001000, 6'b000101, 6'b111000, 6'b100010, 6'b000111, 6'b000000, 6'b000010}, 
{6'b111110, 6'b000010, 6'b000010, 6'b111111, 6'b111101, 6'b111111, 6'b111100, 6'b111111, 6'b000001, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b111110, 6'b111111, 6'b111111, 6'b000010, 6'b111111, 6'b111010, 6'b000011, 6'b000100, 6'b000011, 6'b111101, 6'b111110, 6'b111101, 6'b111101, 6'b000001, 6'b000001, 6'b000001, 6'b000010, 6'b000000, 6'b000011, 6'b111111, 6'b000000, 6'b000010, 6'b000001, 6'b111111, 6'b111111, 6'b000000, 6'b111101, 6'b111110, 6'b111111, 6'b111101, 6'b000011, 6'b000000, 6'b111111, 6'b111111, 6'b111110, 6'b111001, 6'b111111, 6'b111110, 6'b111110, 6'b111111, 6'b000010, 6'b000101, 6'b000001, 6'b111111, 6'b111101, 6'b111111, 6'b000000, 6'b000010, 6'b111111, 6'b000000, 6'b000000}
};

localparam logic signed [5:0] bias [64] = '{
6'b111111,  // -0.037350185215473175
6'b000010,  // 0.27355897426605225
6'b111111,  // -0.12378914654254913
6'b111111,  // -0.064457006752491
6'b000000,  // 0.05452875792980194
6'b000000,  // 0.11671770364046097
6'b000001,  // 0.13640816509723663
6'b000000,  // 0.07482525706291199
6'b000000,  // 0.04674031585454941
6'b111110,  // -0.20146161317825317
6'b111111,  // -0.09910125285387039
6'b000001,  // 0.15104414522647858
6'b111111,  // -0.10221704095602036
6'b111110,  // -0.1461549550294876
6'b111111,  // -0.08641516417264938
6'b000001,  // 0.16613510251045227
6'b111111,  // -0.0836295336484909
6'b111111,  // -0.05756539851427078
6'b111111,  // -0.03229188174009323
6'b111111,  // -0.028388574719429016
6'b000001,  // 0.1260243058204651
6'b111111,  // -0.037064336240291595
6'b000001,  // 0.19336333870887756
6'b000000,  // 0.02124214917421341
6'b000011,  // 0.4985624849796295
6'b000000,  // 0.0158411655575037
6'b111111,  // -0.08296407759189606
6'b000000,  // 0.11056788265705109
6'b000000,  // 0.01173810102045536
6'b111111,  // -0.10843746364116669
6'b000010,  // 0.27439257502555847
6'b000000,  // 0.09199801832437515
6'b000010,  // 0.27419957518577576
6'b000010,  // 0.27063727378845215
6'b111110,  // -0.24828937649726868
6'b000000,  // 0.07818280160427094
6'b111111,  // -0.005749030504375696
6'b000000,  // 0.10850494354963303
6'b000001,  // 0.13591453433036804
6'b111111,  // -0.12088628858327866
6'b111111,  // -0.05666546896100044
6'b000000,  // 0.09311636537313461
6'b000000,  // 0.05477767437696457
6'b000000,  // 0.029585206881165504
6'b111101,  // -0.31209176778793335
6'b111111,  // -0.08465463668107986
6'b111110,  // -0.16775836050510406
6'b000001,  // 0.14762157201766968
6'b111110,  // -0.23618532717227936
6'b000000,  // 0.06535740196704865
6'b111110,  // -0.12853026390075684
6'b111110,  // -0.13802281022071838
6'b111110,  // -0.15156887471675873
6'b000000,  // 0.07979883998632431
6'b000001,  // 0.18141601979732513
6'b111111,  // -0.054039113223552704
6'b111111,  // -0.010052933357656002
6'b000000,  // 0.06611225008964539
6'b000000,  // 0.05053366720676422
6'b000000,  // 0.026860840618610382
6'b000000,  // 0.03283466026186943
6'b000001,  // 0.15558314323425293
6'b111101,  // -0.2863388657569885
6'b111111   // -0.08769102394580841
};
endpackage