// Width: 16
// NFRAC: 6
package dense_3_16_6;

localparam logic signed [15:0] weights [32][32] = '{ 
{16'b1111111111111100, 16'b1111111111100100, 16'b1111111111100110, 16'b1111111111110011, 16'b0000000000010101, 16'b0000000000000010, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000001000, 16'b1111111111011110, 16'b1111111111111100, 16'b0000000000110110, 16'b1111111111110000, 16'b1111111111000100, 16'b1111111111111101, 16'b0000000000000111, 16'b0000000000011011, 16'b1111111111101001, 16'b1111111110111011, 16'b1111111111111101, 16'b0000000000000011, 16'b1111111111100110, 16'b0000000000000000, 16'b0000000001000000, 16'b1111111110100010, 16'b1111111111110001, 16'b1111111111100111, 16'b1111111111110110, 16'b0000000000011011, 16'b1111111111110101}, 
{16'b0000000000101111, 16'b0000000001101110, 16'b0000000000011001, 16'b1111111111010101, 16'b0000000000001111, 16'b1111111111101110, 16'b1111111111111001, 16'b0000000001000101, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111101, 16'b1111111111011010, 16'b1111111111110011, 16'b0000000000100010, 16'b1111111101111001, 16'b1111111111100001, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111100, 16'b1111111111110101, 16'b1111111111101111, 16'b1111111111101110, 16'b0000000000000001, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111110111011, 16'b0000000000000000, 16'b0000000000011110, 16'b1111111111111011, 16'b1111111111010011, 16'b0000000000000000, 16'b0000000000000010}, 
{16'b1111111111000000, 16'b0000000000001011, 16'b0000000000000000, 16'b0000000000010100, 16'b1111111111010111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111001010, 16'b0000000000100010, 16'b1111111111101111, 16'b1111111111101111, 16'b1111111110100000, 16'b1111111111101100, 16'b0000000000100000, 16'b0000000000010000, 16'b1111111111111111, 16'b1111111111111000, 16'b1111111111111110, 16'b1111111111001011, 16'b0000000000000000, 16'b0000000000000111, 16'b0000000000000100, 16'b0000000000001101, 16'b0000000000111000, 16'b0000000000000010, 16'b1111111111001101, 16'b0000000000110001, 16'b0000000000000000, 16'b0000000000001010, 16'b1111111111111110, 16'b0000000000000000, 16'b0000000010010001}, 
{16'b0000000000110101, 16'b1111111111111111, 16'b1111111111110011, 16'b0000000001010011, 16'b0000000001001110, 16'b0000000000000000, 16'b0000000000000100, 16'b0000000000110100, 16'b1111111111100110, 16'b1111111111111111, 16'b1111111111001011, 16'b0000000000000111, 16'b0000000000010001, 16'b1111111111010000, 16'b0000000000000101, 16'b1111111111110101, 16'b1111111111111111, 16'b1111111111101000, 16'b0000000000000010, 16'b0000000000000011, 16'b0000000000000001, 16'b1111111111111011, 16'b0000000001001100, 16'b0000000000101011, 16'b0000000000101010, 16'b0000000000011111, 16'b0000000000101011, 16'b0000000000000000, 16'b1111111111111000, 16'b0000000000111001, 16'b0000000000011111, 16'b1111111111110100}, 
{16'b0000000001000000, 16'b1111111111111010, 16'b1111111111010011, 16'b1111111110011111, 16'b0000000000111101, 16'b0000000000000000, 16'b1111111111001011, 16'b1111111111011011, 16'b1111111111111010, 16'b1111111110011000, 16'b1111111101110010, 16'b0000000000111100, 16'b0000000001010101, 16'b0000000001000010, 16'b1111111110110110, 16'b1111111110011100, 16'b0000000000000000, 16'b1111111111101101, 16'b0000000000011001, 16'b0000000000010001, 16'b1111111111100111, 16'b1111111111111111, 16'b0000000001011100, 16'b1111111101010000, 16'b0000000000001011, 16'b1111111110101011, 16'b0000000000001000, 16'b1111111111100000, 16'b1111111111011001, 16'b1111111111111111, 16'b0000000000001000, 16'b0000000001001010}, 
{16'b0000000000000101, 16'b1111111111111010, 16'b1111111111011000, 16'b1111111111011110, 16'b0000000000101111, 16'b0000000000000000, 16'b1111111111011100, 16'b1111111111101110, 16'b1111111111001001, 16'b1111111111110111, 16'b1111111111111111, 16'b0000000000010100, 16'b0000000000000000, 16'b0000000000101101, 16'b1111111110111111, 16'b1111111111101111, 16'b0000000000001011, 16'b1111111111011010, 16'b1111111111100110, 16'b1111111111111111, 16'b0000000000000001, 16'b0000000000100110, 16'b0000000000111011, 16'b1111111111111110, 16'b1111111111111111, 16'b0000000000110011, 16'b1111111110111001, 16'b1111111111111111, 16'b1111111111100001, 16'b1111111111111011, 16'b1111111111111111, 16'b0000000000000000}, 
{16'b0000000000001000, 16'b1111111111010101, 16'b0000000000001101, 16'b1111111111111011, 16'b1111111111111111, 16'b0000000000010011, 16'b1111111111110010, 16'b1111111110101001, 16'b1111111111111111, 16'b1111111111100101, 16'b1111111111000101, 16'b0000000000111100, 16'b0000000000000000, 16'b0000000001010111, 16'b0000000001101010, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111010111, 16'b1111111111111000, 16'b0000000000100010, 16'b1111111110011111, 16'b0000000000010011, 16'b0000000000101001, 16'b0000000000000010, 16'b0000000000010011, 16'b0000000010011111, 16'b1111111111001101, 16'b1111111111110100, 16'b1111111111100111, 16'b0000000000111110, 16'b1111111111111001, 16'b1111111111101010}, 
{16'b1111111110110011, 16'b0000000000000011, 16'b1111111110101111, 16'b0000000000110111, 16'b0000000010000011, 16'b0000000000001110, 16'b0000000000000000, 16'b0000000000000110, 16'b1111111111111111, 16'b0000000000010000, 16'b0000000010100110, 16'b1111111111111111, 16'b0000000000110000, 16'b0000000001001111, 16'b0000000001100010, 16'b0000000010000110, 16'b0000000000000000, 16'b1111111111000010, 16'b0000000000101011, 16'b1111111111111111, 16'b1111111110101110, 16'b1111111111100010, 16'b0000000000000001, 16'b1111111111110101, 16'b1111111110111111, 16'b0000000011110000, 16'b1111111111100011, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000001110001, 16'b0000000000001011, 16'b0000000000110010}, 
{16'b0000000000110110, 16'b1111111111111101, 16'b0000000000000000, 16'b1111111111111010, 16'b0000000000001010, 16'b1111111111111011, 16'b1111111111111111, 16'b0000000000010100, 16'b0000000000011011, 16'b1111111111011100, 16'b0000000000010001, 16'b0000000000010111, 16'b0000000000000001, 16'b0000000000101010, 16'b1111111111100011, 16'b1111111110011001, 16'b0000000000000000, 16'b1111111111111110, 16'b1111111111111100, 16'b1111111111000000, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111100110, 16'b1111111111111110, 16'b1111111111110011, 16'b0000000000010011, 16'b0000000000101111, 16'b1111111111110000, 16'b1111111111111001, 16'b1111111111111010, 16'b0000000000000011, 16'b1111111111001101}, 
{16'b1111111111101001, 16'b0000000000110001, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000001100101, 16'b0000000000101001, 16'b1111111111111111, 16'b1111111110111000, 16'b0000000000001111, 16'b1111111110100110, 16'b1111111101001100, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000110110, 16'b0000000000001110, 16'b0000000000000000, 16'b1111111111010101, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000111, 16'b0000000000011111, 16'b1111111111111100, 16'b1111111111010001, 16'b0000000000000001, 16'b1111111111111110, 16'b0000000010001010, 16'b0000000000101001, 16'b1111111111111111, 16'b1111111111110110, 16'b0000000001010101, 16'b1111111111111010, 16'b1111111111110100}, 
{16'b1111111110111101, 16'b0000000000010110, 16'b1111111111111011, 16'b1111111111111111, 16'b1111111111100000, 16'b1111111111001111, 16'b0000000000000110, 16'b0000000000010010, 16'b1111111111111111, 16'b1111111111101010, 16'b1111111110110110, 16'b0000000000011001, 16'b0000000000100110, 16'b0000000000000000, 16'b0000000001101011, 16'b1111111110111000, 16'b0000000000001101, 16'b1111111111001101, 16'b0000000000100100, 16'b1111111111111111, 16'b1111111111111011, 16'b0000000000001000, 16'b0000000000001111, 16'b0000000000000000, 16'b1111111111000000, 16'b0000000000000011, 16'b1111111110111000, 16'b1111111111111010, 16'b1111111111111111, 16'b0000000001010110, 16'b1111111111100111, 16'b0000000000000000}, 
{16'b1111111111111111, 16'b0000000000001110, 16'b0000000000000000, 16'b0000000000110010, 16'b1111111111110001, 16'b1111111111111010, 16'b0000000000000111, 16'b1111111111111111, 16'b1111111111111010, 16'b0000000001010010, 16'b0000000001011001, 16'b0000000000000000, 16'b1111111111010101, 16'b1111111110100110, 16'b1111111111111001, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111110111, 16'b1111111111000011, 16'b0000000000110000, 16'b0000000000000000, 16'b0000000000101111, 16'b1111111111111111, 16'b0000000001000111, 16'b0000000000001111, 16'b0000000000100111, 16'b0000000000111010, 16'b1111111111111001, 16'b1111111111001101, 16'b1111111111000111, 16'b1111111111111111, 16'b1111111110101010}, 
{16'b1111111111100011, 16'b1111111111111111, 16'b0000000000001111, 16'b1111111111001010, 16'b0000000000001011, 16'b1111111111111111, 16'b1111111111100100, 16'b1111111111111110, 16'b1111111111101111, 16'b0000000000000100, 16'b0000000000001001, 16'b1111111111110110, 16'b0000000000000010, 16'b0000000000011000, 16'b1111111110101111, 16'b1111111111100000, 16'b0000000000011101, 16'b1111111111101001, 16'b0000000000000000, 16'b1111111111111100, 16'b0000000000011000, 16'b0000000000000001, 16'b1111111111111100, 16'b0000000000000101, 16'b0000000000100010, 16'b1111111111110010, 16'b0000000000000000, 16'b1111111111000110, 16'b1111111111100110, 16'b1111111111111111, 16'b0000000000010110, 16'b0000000000000000}, 
{16'b1111111110111101, 16'b0000000000110101, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111110, 16'b0000000000010110, 16'b1111111111111111, 16'b0000000001100010, 16'b1111111111111110, 16'b1111111111111111, 16'b0000000000011010, 16'b0000000000000101, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000001111, 16'b0000000000101010, 16'b0000000000010110, 16'b0000000000010101, 16'b1111111111111110, 16'b0000000000100111, 16'b0000000000001100, 16'b0000000000000101, 16'b1111111111111110, 16'b0000000000100000, 16'b1111111111110011, 16'b1111111111010100, 16'b1111111111110100, 16'b1111111111111111, 16'b0000000000001101, 16'b0000000000000011, 16'b0000000000011001, 16'b0000000000111101}, 
{16'b1111111111111101, 16'b1111111111001110, 16'b0000000000000110, 16'b1111111111111111, 16'b0000000001110101, 16'b1111111111100101, 16'b1111111110110110, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111100, 16'b0000000000000110, 16'b0000000000110111, 16'b0000000000101001, 16'b0000000000000001, 16'b0000000000000100, 16'b1111111111101001, 16'b0000000000000100, 16'b1111111111111011, 16'b0000000000000000, 16'b0000000000001001, 16'b1111111111111011, 16'b0000000000000010, 16'b0000000000100010, 16'b0000000000000100, 16'b1111111111111110, 16'b1111111111001011, 16'b0000000000011010, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111110010, 16'b1111111111111101, 16'b1111111111110111}, 
{16'b0000000000000000, 16'b1111111111110111, 16'b1111111111101111, 16'b1111111111100100, 16'b1111111110111010, 16'b0000000001001110, 16'b0000000000000000, 16'b0000000000010101, 16'b0000000000100100, 16'b0000000000000001, 16'b1111111111111011, 16'b0000000000111100, 16'b0000000000011100, 16'b1111111111010001, 16'b1111111111101011, 16'b1111111111111010, 16'b1111111111001101, 16'b1111111111111101, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000010011, 16'b1111111111101110, 16'b0000000000000000, 16'b0000000000001001, 16'b1111111111111111, 16'b1111111111010100, 16'b0000000000010100, 16'b0000000000000000, 16'b0000000000000101, 16'b0000000000000001, 16'b1111111111010111, 16'b0000000000000010}, 
{16'b1111111111100110, 16'b1111111111101011, 16'b0000000000001001, 16'b1111111111110000, 16'b1111111111110100, 16'b0000000000001110, 16'b1111111111111111, 16'b0000000000000100, 16'b0000000000010000, 16'b1111111111111111, 16'b0000000000001111, 16'b1111111111101111, 16'b1111111111111110, 16'b1111111111111111, 16'b0000000000001101, 16'b1111111111111111, 16'b0000000000111110, 16'b1111111111111101, 16'b0000000000011111, 16'b1111111111101010, 16'b0000000000010100, 16'b0000000000001000, 16'b0000000000001010, 16'b0000000000000100, 16'b1111111111110101, 16'b1111111111011100, 16'b1111111111011110, 16'b0000000000001101, 16'b1111111111110101, 16'b0000000000000000, 16'b1111111111111100, 16'b0000000000011101}, 
{16'b1111111111111111, 16'b1111111111001100, 16'b1111111111001101, 16'b1111111111111111, 16'b0000000001010000, 16'b1111111111110100, 16'b0000000000000000, 16'b0000000000111101, 16'b1111111111101101, 16'b0000000000000000, 16'b1111111111001010, 16'b1111111111000001, 16'b0000000000111001, 16'b0000000000010011, 16'b1111111111110000, 16'b1111111111011100, 16'b0000000000010110, 16'b0000000000000000, 16'b1111111111100001, 16'b0000000000000011, 16'b0000000000001000, 16'b1111111111110100, 16'b0000000000100100, 16'b1111111110000010, 16'b0000000000000101, 16'b0000000000011110, 16'b1111111111111010, 16'b0000000000000001, 16'b1111111111100010, 16'b1111111111111111, 16'b1111111111100110, 16'b1111111111111100}, 
{16'b0000000000011011, 16'b0000000000101100, 16'b0000000001000110, 16'b1111111111100101, 16'b0000000000110101, 16'b0000000000100111, 16'b0000000000000000, 16'b0000000000111010, 16'b0000000000101101, 16'b1111111111110010, 16'b0000000001011001, 16'b1111111111010011, 16'b0000000001001111, 16'b0000000000111001, 16'b1111111101110110, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000100001, 16'b1111111110111111, 16'b0000000000011100, 16'b1111111111100100, 16'b1111111111000001, 16'b1111111111101011, 16'b0000000000101010, 16'b1111111110101011, 16'b1111111111010101, 16'b1111111111111010, 16'b1111111111111111, 16'b1111111110110111, 16'b0000000000110010, 16'b0000000000000000}, 
{16'b1111111111111001, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111010011, 16'b0000000000000001, 16'b0000000000000001, 16'b1111111111111110, 16'b1111111111111100, 16'b1111111111111010, 16'b0000000000010001, 16'b1111111111111111, 16'b0000000000001010, 16'b1111111111010100, 16'b0000000000001101, 16'b1111111111111111, 16'b0000000000010010, 16'b0000000000111001, 16'b1111111111010010, 16'b0000000000000110, 16'b1111111111110011, 16'b0000000000010000, 16'b0000000000011000, 16'b1111111111110101, 16'b1111111111011111, 16'b0000000000000010, 16'b0000000001101010, 16'b1111111111111100, 16'b1111111111111110, 16'b0000000000101001, 16'b0000000000000000, 16'b0000000001101110}, 
{16'b1111111110111101, 16'b0000000000000100, 16'b1111111111100100, 16'b0000000000110001, 16'b0000000000001110, 16'b1111111111111011, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111011001, 16'b1111111111111011, 16'b0000000000000000, 16'b1111111110111000, 16'b0000000000000001, 16'b1111111111111010, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111110001, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000010100, 16'b0000000000000010, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111110, 16'b0000000000000000, 16'b0000000000000010, 16'b0000000001001010, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111010, 16'b0000000000010110, 16'b1111111111111100}, 
{16'b1111111111111111, 16'b1111111111101100, 16'b0000000000011010, 16'b0000000000000101, 16'b1111111111010000, 16'b0000000000000000, 16'b0000000000100100, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111110011, 16'b0000000000001110, 16'b0000000000000010, 16'b0000000000101001, 16'b1111111110111001, 16'b1111111111110011, 16'b1111111111111101, 16'b0000000000011011, 16'b1111111111001110, 16'b0000000000000010, 16'b1111111110011111, 16'b1111111111111101, 16'b1111111111110000, 16'b1111111111111010, 16'b0000000000100101, 16'b1111111111110110, 16'b1111111111011100, 16'b0000000000001011, 16'b0000000000000000, 16'b0000000000110010, 16'b0000000001000010, 16'b1111111111010110, 16'b1111111111000110}, 
{16'b0000000000001000, 16'b0000000000000011, 16'b1111111111001010, 16'b1111111111111000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000001101, 16'b0000000000110100, 16'b0000000000000000, 16'b0000000000000010, 16'b0000000000001000, 16'b1111111110111010, 16'b1111111111110111, 16'b1111111110110010, 16'b0000000000111101, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111110101101, 16'b1111111111111111, 16'b1111111111110110, 16'b1111111111111101, 16'b0000000000000000, 16'b0000000000000111, 16'b1111111111101100, 16'b0000000000000110, 16'b0000000000110100, 16'b0000000000110110, 16'b0000000000110001, 16'b0000000000100111, 16'b0000000000000000, 16'b0000000000001110, 16'b0000000001100100}, 
{16'b1111111111111100, 16'b1111111111100001, 16'b0000000000110001, 16'b1111111111110010, 16'b0000000000001000, 16'b0000000000010101, 16'b1111111111111111, 16'b1111111111011011, 16'b1111111111110101, 16'b1111111110110011, 16'b0000000000111001, 16'b0000000000000000, 16'b0000000000110101, 16'b0000000001010101, 16'b1111111111110001, 16'b1111111110010000, 16'b1111111111110010, 16'b0000000000111100, 16'b1111111111011011, 16'b1111111111100101, 16'b0000000000000111, 16'b0000000000000000, 16'b1111111110111010, 16'b1111111111100111, 16'b1111111111111010, 16'b1111111111110000, 16'b0000000000001110, 16'b0000000001011010, 16'b0000000000011111, 16'b1111111111111111, 16'b0000000000001010, 16'b0000000000000011}, 
{16'b0000000000000101, 16'b0000000000111010, 16'b0000000000000000, 16'b0000000000100101, 16'b0000000001101010, 16'b1111111111101010, 16'b1111111111111111, 16'b1111111111111010, 16'b0000000000100101, 16'b1111111111100111, 16'b1111111111111111, 16'b0000000000101010, 16'b0000000000000001, 16'b0000000000000011, 16'b1111111100111100, 16'b1111111111110101, 16'b0000000000000000, 16'b0000000000011001, 16'b1111111111111111, 16'b0000000000100110, 16'b1111111111111111, 16'b1111111111101001, 16'b1111111110111000, 16'b0000000000010000, 16'b0000000000100100, 16'b1111111101110010, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000001000101, 16'b1111111110011001, 16'b0000000000000000, 16'b1111111111111111}, 
{16'b0000000000000001, 16'b1111111111010100, 16'b0000000000000110, 16'b1111111111111110, 16'b0000000000000110, 16'b0000000001000011, 16'b1111111110100011, 16'b0000000000000100, 16'b0000000000110110, 16'b1111111111010100, 16'b1111111111111101, 16'b0000000000000110, 16'b1111111111111110, 16'b0000000000010110, 16'b0000000000001101, 16'b1111111111111101, 16'b0000000000001000, 16'b0000000000000000, 16'b0000000000000010, 16'b0000000000110000, 16'b1111111111111100, 16'b1111111111000010, 16'b1111111110110010, 16'b1111111111100111, 16'b1111111110110100, 16'b0000000000011010, 16'b0000000001001111, 16'b0000000000101111, 16'b1111111111111110, 16'b1111111111010000, 16'b1111111111011000, 16'b0000000000000111}, 
{16'b0000000000000110, 16'b1111111111000010, 16'b1111111111111101, 16'b0000000000010011, 16'b1111111111000010, 16'b0000000000010101, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000100001, 16'b1111111111111101, 16'b0000000000000001, 16'b0000000000000000, 16'b0000000000010000, 16'b1111111111111101, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111010110, 16'b1111111110111111, 16'b1111111111111111, 16'b1111111110111011, 16'b1111111111011001, 16'b1111111111010000, 16'b0000000001110001, 16'b0000000000000010, 16'b1111111111111010, 16'b0000000000101000, 16'b0000000001110010, 16'b0000000000110010, 16'b1111111101111000, 16'b1111111111101000}, 
{16'b0000000000110000, 16'b1111111111111111, 16'b0000000000100000, 16'b1111111111111101, 16'b0000000000111101, 16'b1111111111101101, 16'b0000000000001001, 16'b0000000000110101, 16'b0000000000100010, 16'b1111111110111101, 16'b1111111111111000, 16'b0000000000001111, 16'b0000000000001000, 16'b1111111111111110, 16'b0000000000001010, 16'b0000000000000000, 16'b0000000000101110, 16'b0000000000000100, 16'b0000000000101111, 16'b1111111111110111, 16'b1111111111101111, 16'b1111111111110110, 16'b1111111111111111, 16'b0000000000100110, 16'b1111111111100110, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000100101, 16'b1111111111010110, 16'b1111111111111101}, 
{16'b1111111111111111, 16'b1111111111111100, 16'b1111111111000100, 16'b0000000000100100, 16'b0000000000011100, 16'b1111111111110001, 16'b1111111111111111, 16'b1111111111100010, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111011001, 16'b1111111111100000, 16'b0000000000111101, 16'b0000000000000000, 16'b1111111111101111, 16'b1111111111111111, 16'b0000000000011011, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111100100, 16'b0000000000101000, 16'b0000000000000000, 16'b0000000000010011, 16'b1111111111111100, 16'b0000000000010100, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000011110, 16'b1111111111100111, 16'b1111111111111010, 16'b0000000000010100, 16'b1111111111110010}, 
{16'b1111111111111101, 16'b1111111111011000, 16'b0000000001001100, 16'b1111111111110111, 16'b0000000000011001, 16'b1111111111011011, 16'b0000000000000000, 16'b0000000000000100, 16'b1111111111000010, 16'b1111111111111110, 16'b1111111111110000, 16'b0000000000000111, 16'b1111111111010110, 16'b0000000000010001, 16'b0000000000011001, 16'b0000000000001110, 16'b0000000000001010, 16'b1111111111111011, 16'b1111111110100101, 16'b1111111111111110, 16'b1111111111111000, 16'b0000000000010001, 16'b1111111111110001, 16'b1111111111111111, 16'b0000000000011001, 16'b1111111111111010, 16'b1111111111111110, 16'b0000000000110001, 16'b1111111111001101, 16'b1111111111011010, 16'b0000000000101100, 16'b0000000000000100}, 
{16'b0000000000110111, 16'b0000000000011001, 16'b0000000000000000, 16'b1111111111101011, 16'b1111111111110101, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111110111, 16'b1111111111110000, 16'b1111111111110000, 16'b0000000000000000, 16'b0000000000010100, 16'b0000000000000000, 16'b0000000000000110, 16'b1111111111111010, 16'b0000000000000000, 16'b1111111111101100, 16'b0000000000000000, 16'b1111111111111101, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000111, 16'b0000000000001100, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111110110001, 16'b1111111111100110, 16'b0000000000000000, 16'b0000000000000010, 16'b0000000000000000, 16'b1111111111101001, 16'b0000000000000010}, 
{16'b0000000000011000, 16'b1111111101111010, 16'b1111111111111111, 16'b1111111111110110, 16'b1111111111100010, 16'b1111111111111110, 16'b0000000000000000, 16'b0000000001000110, 16'b1111111111111010, 16'b1111111111111101, 16'b0000000000001010, 16'b1111111110101011, 16'b0000000000000011, 16'b1111111111000111, 16'b0000000001011100, 16'b1111111111111001, 16'b1111111111100011, 16'b1111111110111001, 16'b1111111111111110, 16'b1111111110100101, 16'b1111111110011000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000011111, 16'b1111111111111110, 16'b1111111111011001, 16'b1111111111110110, 16'b1111111111111101, 16'b0000000000000000, 16'b1111111111111011, 16'b1111111110100110}
};

localparam logic signed [15:0] bias [32] = '{
16'b0000000000100001,  // 0.5280959606170654
16'b0000000000110101,  // 0.8414360880851746
16'b0000000000011001,  // 0.397830605506897
16'b0000000000011010,  // 0.4105983078479767
16'b1111111100010101,  // -3.657735586166382
16'b1111111111000110,  // -0.8977976441383362
16'b0000000001101101,  // 1.7051936388015747
16'b1111111110101110,  // -1.2765135765075684
16'b1111111111011010,  // -0.5837795734405518
16'b0000000010101100,  // 2.699671983718872
16'b0000000000001101,  // 0.2170683741569519
16'b0000000000111000,  // 0.8814588785171509
16'b1111111101010111,  // -2.634300947189331
16'b1111111110000111,  // -1.877297282218933
16'b0000000001101010,  // 1.6625694036483765
16'b0000000010101111,  // 2.7459704875946045
16'b1111111111100001,  // -0.47838035225868225
16'b0000000001101100,  // 1.6984987258911133
16'b0000000000110110,  // 0.8548859357833862
16'b0000000001000000,  // 1.0045719146728516
16'b0000000001011010,  // 1.4197649955749512
16'b0000000000110101,  // 0.832463800907135
16'b0000000000100010,  // 0.5434179306030273
16'b0000000000111011,  // 0.9277304410934448
16'b1111111111101010,  // -0.3426123857498169
16'b1111111111011100,  // -0.5587119460105896
16'b1111111111011000,  // -0.6208624839782715
16'b1111111110101110,  // -1.2802538871765137
16'b0000000000000011,  // 0.05940237268805504
16'b1111111111001011,  // -0.8213341236114502
16'b0000000000111000,  // 0.8783953189849854
16'b1111111111000011   // -0.949700653553009
};
endpackage