// Width: 23
// NFRAC: 11
package dense_4_23_11;

localparam logic signed [22:0] weights [32][5] = '{ 
{23'b11111111111111111100111, 23'b00000000000001010000110, 23'b11111111111110110011101, 23'b00000000000000010000110, 23'b11111111111111100100110}, 
{23'b11111111111101110001001, 23'b11111111111111110001111, 23'b00000000000001110101110, 23'b11111111111111111100110, 23'b00000000000000000100010}, 
{23'b00000000000001011111000, 23'b00000000000000110110001, 23'b11111111111111111000110, 23'b11111111111110011000001, 23'b11111111111111001010000}, 
{23'b11111111111110011111110, 23'b11111111111110100000100, 23'b11111111111111100011011, 23'b00000000000001001110110, 23'b00000000000000111100001}, 
{23'b00000000000000011111010, 23'b00000000000000100000111, 23'b00000000000000101000001, 23'b11111111111111111011010, 23'b11111111111011111100101}, 
{23'b00000000000001010011101, 23'b11111111111110011011000, 23'b00000000000000101110011, 23'b11111111111111010110101, 23'b11111111111111010100011}, 
{23'b11111111111110011001010, 23'b00000000000000001001000, 23'b11111111111111111111111, 23'b00000000000000101100100, 23'b00000000000000010001101}, 
{23'b11111111111111111111100, 23'b00000000000001001000110, 23'b11111111111110011011101, 23'b00000000000000101001101, 23'b00000000000000100010110}, 
{23'b00000000000000101001110, 23'b11111111111111010100101, 23'b00000000000000000000010, 23'b11111111111110001001110, 23'b11111111111111000000010}, 
{23'b11111111111111111111111, 23'b11111111111110111011110, 23'b00000000000000101101100, 23'b00000000000001101110000, 23'b00000000000000000000000}, 
{23'b11111111111111011110101, 23'b11111111111111011010111, 23'b00000000000000000000000, 23'b00000000000010010100110, 23'b11111111111110111011011}, 
{23'b00000000000000101011010, 23'b00000000000000111010101, 23'b11111111111110101000111, 23'b11111111111111111000111, 23'b00000000000000011111001}, 
{23'b00000000000000000000000, 23'b00000000000000101010111, 23'b00000000000000000010010, 23'b11111111111111001010110, 23'b11111111111101100000100}, 
{23'b00000000000000101101011, 23'b00000000000000010000010, 23'b00000000000001101011011, 23'b11111111111111101110000, 23'b11111111111110010010011}, 
{23'b00000000000000010111001, 23'b11111111111111110011101, 23'b11111111111110100011101, 23'b11111111111111110111100, 23'b00000000000010001001010}, 
{23'b11111111111110000110101, 23'b11111111111111000001011, 23'b11111111111111000111000, 23'b00000000000001100110000, 23'b00000000000000001000001}, 
{23'b00000000000001011000100, 23'b11111111111111010100000, 23'b11111111111111011101010, 23'b11111111111111000110001, 23'b11111111111111110000101}, 
{23'b00000000000000110001111, 23'b11111111111111110101101, 23'b11111111111110010110011, 23'b11111111111111111000001, 23'b00000000000000010010000}, 
{23'b00000000000001000010001, 23'b00000000000000001010101, 23'b11111111111111001000001, 23'b00000000000000000000000, 23'b11111111111110011111110}, 
{23'b00000000000000111011001, 23'b11111111111111101001110, 23'b11111111111111001001100, 23'b00000000000000110101000, 23'b00000000000000011000010}, 
{23'b00000000000000010001010, 23'b11111111111111111000001, 23'b00000000000001001100001, 23'b11111111111110010001101, 23'b11111111111111111010100}, 
{23'b00000000000000000000000, 23'b00000000000000011110001, 23'b00000000000001111100100, 23'b11111111111101111011010, 23'b11111111111101100001111}, 
{23'b11111111111111100110110, 23'b00000000000000011100000, 23'b00000000000000101101010, 23'b11111111111110100100101, 23'b00000000000010000101101}, 
{23'b11111111111111111111111, 23'b00000000000000101010001, 23'b00000000000001001000010, 23'b00000000000000001001101, 23'b11111111111101101101100}, 
{23'b11111111111111010100101, 23'b00000000000001011101010, 23'b11111111111111000110110, 23'b00000000000000000001011, 23'b00000000000001100011010}, 
{23'b00000000000000000110101, 23'b00000000000001000100000, 23'b00000000000000000111100, 23'b11111111111101000000100, 23'b00000000000010001100010}, 
{23'b11111111111110001010010, 23'b11111111111111000001101, 23'b00000000000000110110110, 23'b00000000000000111110100, 23'b00000000000000110011101}, 
{23'b00000000000000000001000, 23'b00000000000000111101101, 23'b11111111111111110110101, 23'b11111111111111011001011, 23'b00000000000000001000000}, 
{23'b11111111111111100101010, 23'b00000000000000111111000, 23'b11111111111101111111000, 23'b00000000000000100011100, 23'b11111111111111010111011}, 
{23'b11111111111111111011010, 23'b00000000000000100100001, 23'b11111111111111010100110, 23'b11111111111110011001011, 23'b00000000000010010111111}, 
{23'b00000000000001110010111, 23'b00000000000000010001111, 23'b00000000000001010011000, 23'b11111111111101101001000, 23'b11111111111110101111010}, 
{23'b11111111111111110000110, 23'b11111111111110011101001, 23'b00000000000001011101101, 23'b00000000000000010010001, 23'b00000000000000100000101}
};

localparam logic signed [22:0] bias [5] = '{
23'b11111111111111110000000,  // -0.06223141402006149
23'b11111111111111101111111,  // -0.06270556896924973
23'b11111111111111101110000,  // -0.07014333456754684
23'b00000000000000010101000,  // 0.0820775106549263
23'b00000000000000110111001   // 0.2155742198228836
};
endpackage