// Width: 18
// NFRAC: 9
package dense_3_18_9;

localparam logic signed [17:0] weights [32][32] = '{ 
{18'b111111111111100110, 18'b111111111100100000, 18'b111111111100110000, 18'b111111111110011110, 18'b000000000010101111, 18'b000000000000010110, 18'b111111111111111001, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000001000000, 18'b111111111011110010, 18'b111111111111100001, 18'b000000000110110001, 18'b111111111110000100, 18'b111111111000100010, 18'b111111111111101101, 18'b000000000000111001, 18'b000000000011011110, 18'b111111111101001101, 18'b111111110111011110, 18'b111111111111101000, 18'b000000000000011001, 18'b111111111100110001, 18'b000000000000000000, 18'b000000001000000110, 18'b111111110100010110, 18'b111111111110001110, 18'b111111111100111001, 18'b111111111110110011, 18'b000000000011011000, 18'b111111111110101110}, 
{18'b000000000101111110, 18'b000000001101110101, 18'b000000000011001101, 18'b111111111010101111, 18'b000000000001111101, 18'b111111111101110100, 18'b111111111111001000, 18'b000000001000101110, 18'b000000000000000011, 18'b111111111111111111, 18'b111111111111101111, 18'b111111111011010010, 18'b111111111110011000, 18'b000000000100010100, 18'b111111101111001001, 18'b111111111100001110, 18'b111111111111111111, 18'b111111111111111011, 18'b111111111111100101, 18'b111111111110101011, 18'b111111111101111011, 18'b111111111101110011, 18'b000000000000001000, 18'b111111111111111111, 18'b111111111111111100, 18'b111111110111011011, 18'b000000000000000110, 18'b000000000011110001, 18'b111111111111011111, 18'b111111111010011110, 18'b000000000000000001, 18'b000000000000010011}, 
{18'b111111111000000111, 18'b000000000001011110, 18'b000000000000000101, 18'b000000000010100101, 18'b111111111010111101, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111001010010, 18'b000000000100010010, 18'b111111111101111001, 18'b111111111101111011, 18'b111111110100000110, 18'b111111111101100000, 18'b000000000100000101, 18'b000000000010000111, 18'b111111111111111111, 18'b111111111111000101, 18'b111111111111110011, 18'b111111111001011110, 18'b000000000000000001, 18'b000000000000111111, 18'b000000000000100011, 18'b000000000001101011, 18'b000000000111000010, 18'b000000000000010011, 18'b111111111001101100, 18'b000000000110001000, 18'b000000000000000000, 18'b000000000001010100, 18'b111111111111110100, 18'b000000000000000000, 18'b000000010010001001}, 
{18'b000000000110101100, 18'b111111111111111111, 18'b111111111110011100, 18'b000000001010011110, 18'b000000001001110100, 18'b000000000000000000, 18'b000000000000100101, 18'b000000000110100000, 18'b111111111100110101, 18'b111111111111111111, 18'b111111111001011010, 18'b000000000000111101, 18'b000000000010001000, 18'b111111111010000001, 18'b000000000000101111, 18'b111111111110101110, 18'b111111111111111111, 18'b111111111101000101, 18'b000000000000010011, 18'b000000000000011100, 18'b000000000000001000, 18'b111111111111011010, 18'b000000001001100011, 18'b000000000101011111, 18'b000000000101010001, 18'b000000000011111110, 18'b000000000101011101, 18'b000000000000000000, 18'b111111111111000011, 18'b000000000111001111, 18'b000000000011111111, 18'b111111111110100110}, 
{18'b000000001000000000, 18'b111111111111010000, 18'b111111111010011101, 18'b111111110011111110, 18'b000000000111101000, 18'b000000000000000000, 18'b111111111001011011, 18'b111111111011011110, 18'b111111111111010000, 18'b111111110011000011, 18'b111111101110010100, 18'b000000000111100100, 18'b000000001010101100, 18'b000000001000010111, 18'b111111110110110011, 18'b111111110011100110, 18'b000000000000000000, 18'b111111111101101111, 18'b000000000011001101, 18'b000000000010001110, 18'b111111111100111111, 18'b111111111111111001, 18'b000000001011100010, 18'b111111101010000000, 18'b000000000001011010, 18'b111111110101011101, 18'b000000000001000011, 18'b111111111100000001, 18'b111111111011001110, 18'b111111111111111111, 18'b000000000001000111, 18'b000000001001010010}, 
{18'b000000000000101100, 18'b111111111111010101, 18'b111111111011000101, 18'b111111111011110101, 18'b000000000101111100, 18'b000000000000000000, 18'b111111111011100001, 18'b111111111101110100, 18'b111111111001001001, 18'b111111111110111110, 18'b111111111111111111, 18'b000000000010100100, 18'b000000000000000000, 18'b000000000101101110, 18'b111111110111111010, 18'b111111111101111101, 18'b000000000001011011, 18'b111111111011010011, 18'b111111111100110101, 18'b111111111111111111, 18'b000000000000001100, 18'b000000000100110010, 18'b000000000111011110, 18'b111111111111110101, 18'b111111111111111111, 18'b000000000110011010, 18'b111111110111001101, 18'b111111111111111111, 18'b111111111100001101, 18'b111111111111011010, 18'b111111111111111100, 18'b000000000000000110}, 
{18'b000000000001000010, 18'b111111111010101011, 18'b000000000001101110, 18'b111111111111011000, 18'b111111111111111000, 18'b000000000010011011, 18'b111111111110010011, 18'b111111110101001010, 18'b111111111111111111, 18'b111111111100101010, 18'b111111111000101100, 18'b000000000111100011, 18'b000000000000000111, 18'b000000001010111100, 18'b000000001101010000, 18'b000000000000000010, 18'b111111111111111111, 18'b111111111010111101, 18'b111111111111000000, 18'b000000000100010111, 18'b111111110011111111, 18'b000000000010011111, 18'b000000000101001110, 18'b000000000000010011, 18'b000000000010011001, 18'b000000010011111001, 18'b111111111001101100, 18'b111111111110100011, 18'b111111111100111101, 18'b000000000111110010, 18'b111111111111001101, 18'b111111111101010010}, 
{18'b111111110110011101, 18'b000000000000011000, 18'b111111110101111011, 18'b000000000110111101, 18'b000000010000011100, 18'b000000000001110110, 18'b000000000000000011, 18'b000000000000110000, 18'b111111111111111111, 18'b000000000010000011, 18'b000000010100110100, 18'b111111111111111111, 18'b000000000110000110, 18'b000000001001111101, 18'b000000001100010011, 18'b000000010000110011, 18'b000000000000000000, 18'b111111111000010110, 18'b000000000101011000, 18'b111111111111111010, 18'b111111110101110010, 18'b111111111100010111, 18'b000000000000001101, 18'b111111111110101011, 18'b111111110111111110, 18'b000000011110000000, 18'b111111111100011111, 18'b000000000000000000, 18'b000000000000000000, 18'b000000001110001000, 18'b000000000001011010, 18'b000000000110010001}, 
{18'b000000000110110000, 18'b111111111111101100, 18'b000000000000000000, 18'b111111111111010011, 18'b000000000001010011, 18'b111111111111011001, 18'b111111111111111111, 18'b000000000010100000, 18'b000000000011011000, 18'b111111111011100111, 18'b000000000010001111, 18'b000000000010111111, 18'b000000000000001100, 18'b000000000101010100, 18'b111111111100011001, 18'b111111110011001111, 18'b000000000000000000, 18'b111111111111110001, 18'b111111111111100100, 18'b111111111000000001, 18'b111111111111111110, 18'b000000000000000000, 18'b111111111100110000, 18'b111111111111110001, 18'b111111111110011110, 18'b000000000010011111, 18'b000000000101111110, 18'b111111111110000101, 18'b111111111111001101, 18'b111111111111010110, 18'b000000000000011011, 18'b111111111001101110}, 
{18'b111111111101001010, 18'b000000000110001001, 18'b000000000000000000, 18'b000000000000000000, 18'b000000001100101011, 18'b000000000101001001, 18'b111111111111111111, 18'b111111110111000111, 18'b000000000001111000, 18'b111111110100110101, 18'b111111101001100011, 18'b111111111111111111, 18'b000000000000000000, 18'b000000000110110111, 18'b000000000001110001, 18'b000000000000000000, 18'b111111111010101111, 18'b000000000000000000, 18'b000000000000000110, 18'b000000000000111110, 18'b000000000011111001, 18'b111111111111100101, 18'b111111111010001111, 18'b000000000000001000, 18'b111111111111110100, 18'b000000010001010011, 18'b000000000101001110, 18'b111111111111111111, 18'b111111111110110111, 18'b000000001010101100, 18'b111111111111010111, 18'b111111111110100110}, 
{18'b111111110111101000, 18'b000000000010110011, 18'b111111111111011100, 18'b111111111111111111, 18'b111111111100000011, 18'b111111111001111101, 18'b000000000000110001, 18'b000000000010010011, 18'b111111111111111111, 18'b111111111101010000, 18'b111111110110110101, 18'b000000000011001101, 18'b000000000100110111, 18'b000000000000000000, 18'b000000001101011011, 18'b111111110111000000, 18'b000000000001101010, 18'b111111111001101111, 18'b000000000100100000, 18'b111111111111111111, 18'b111111111111011000, 18'b000000000001000111, 18'b000000000001111101, 18'b000000000000000000, 18'b111111111000000110, 18'b000000000000011111, 18'b111111110111000011, 18'b111111111111010111, 18'b111111111111111111, 18'b000000001010110011, 18'b111111111100111101, 18'b000000000000000000}, 
{18'b111111111111111111, 18'b000000000001110101, 18'b000000000000000000, 18'b000000000110010000, 18'b111111111110001000, 18'b111111111111010011, 18'b000000000000111011, 18'b111111111111111010, 18'b111111111111010000, 18'b000000001010010000, 18'b000000001011001011, 18'b000000000000000000, 18'b111111111010101011, 18'b111111110100110000, 18'b111111111111001100, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111110111110, 18'b111111111000011000, 18'b000000000110000111, 18'b000000000000000010, 18'b000000000101111011, 18'b111111111111111111, 18'b000000001000111111, 18'b000000000001111110, 18'b000000000100111001, 18'b000000000111010010, 18'b111111111111001011, 18'b111111111001101111, 18'b111111111000111100, 18'b111111111111111010, 18'b111111110101010011}, 
{18'b111111111100011000, 18'b111111111111111111, 18'b000000000001111010, 18'b111111111001010011, 18'b000000000001011000, 18'b111111111111111111, 18'b111111111100100001, 18'b111111111111110110, 18'b111111111101111111, 18'b000000000000100110, 18'b000000000001001111, 18'b111111111110110110, 18'b000000000000010000, 18'b000000000011000000, 18'b111111110101111111, 18'b111111111100000101, 18'b000000000011101001, 18'b111111111101001010, 18'b000000000000000000, 18'b111111111111100110, 18'b000000000011000101, 18'b000000000000001000, 18'b111111111111100000, 18'b000000000000101011, 18'b000000000100010011, 18'b111111111110010101, 18'b000000000000000000, 18'b111111111000110001, 18'b111111111100110111, 18'b111111111111111000, 18'b000000000010110001, 18'b000000000000000000}, 
{18'b111111110111101011, 18'b000000000110101110, 18'b111111111111111111, 18'b111111111111111001, 18'b111111111111110110, 18'b000000000010110011, 18'b111111111111111111, 18'b000000001100010110, 18'b111111111111110000, 18'b111111111111111111, 18'b000000000011010010, 18'b000000000000101001, 18'b000000000000000110, 18'b000000000000000000, 18'b000000000001111100, 18'b000000000101010010, 18'b000000000010110110, 18'b000000000010101010, 18'b111111111111110111, 18'b000000000100111010, 18'b000000000001100111, 18'b000000000000101001, 18'b111111111111110111, 18'b000000000100000100, 18'b111111111110011010, 18'b111111111010100100, 18'b111111111110100001, 18'b111111111111111111, 18'b000000000001101000, 18'b000000000000011110, 18'b000000000011001000, 18'b000000000111101010}, 
{18'b111111111111101100, 18'b111111111001110001, 18'b000000000000110100, 18'b111111111111111111, 18'b000000001110101010, 18'b111111111100101011, 18'b111111110110110110, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111111100101, 18'b000000000000110001, 18'b000000000110111111, 18'b000000000101001001, 18'b000000000000001010, 18'b000000000000100010, 18'b111111111101001101, 18'b000000000000100010, 18'b111111111111011001, 18'b000000000000000000, 18'b000000000001001101, 18'b111111111111011001, 18'b000000000000010011, 18'b000000000100010000, 18'b000000000000100101, 18'b111111111111110011, 18'b111111111001011001, 18'b000000000011010000, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111110010011, 18'b111111111111101010, 18'b111111111110111111}, 
{18'b000000000000000111, 18'b111111111110111111, 18'b111111111101111110, 18'b111111111100100000, 18'b111111110111010000, 18'b000000001001110000, 18'b000000000000000000, 18'b000000000010101100, 18'b000000000100100101, 18'b000000000000001101, 18'b111111111111011101, 18'b000000000111100111, 18'b000000000011100101, 18'b111111111010001001, 18'b111111111101011001, 18'b111111111111010101, 18'b111111111001101000, 18'b111111111111101110, 18'b000000000000000000, 18'b111111111111111011, 18'b000000000010011111, 18'b111111111101110011, 18'b000000000000000000, 18'b000000000001001110, 18'b111111111111111111, 18'b111111111010100010, 18'b000000000010100000, 18'b000000000000000000, 18'b000000000000101101, 18'b000000000000001011, 18'b111111111010111100, 18'b000000000000010101}, 
{18'b111111111100110111, 18'b111111111101011110, 18'b000000000001001110, 18'b111111111110000000, 18'b111111111110100100, 18'b000000000001110110, 18'b111111111111111010, 18'b000000000000100011, 18'b000000000010000110, 18'b111111111111111111, 18'b000000000001111110, 18'b111111111101111101, 18'b111111111111110110, 18'b111111111111111111, 18'b000000000001101001, 18'b111111111111111111, 18'b000000000111110100, 18'b111111111111101110, 18'b000000000011111110, 18'b111111111101010010, 18'b000000000010100010, 18'b000000000001000000, 18'b000000000001010110, 18'b000000000000100101, 18'b111111111110101100, 18'b111111111011100010, 18'b111111111011110110, 18'b000000000001101110, 18'b111111111110101010, 18'b000000000000000000, 18'b111111111111100011, 18'b000000000011101101}, 
{18'b111111111111111111, 18'b111111111001100001, 18'b111111111001101001, 18'b111111111111111111, 18'b000000001010000110, 18'b111111111110100011, 18'b000000000000000000, 18'b000000000111101110, 18'b111111111101101000, 18'b000000000000000000, 18'b111111111001010100, 18'b111111111000001010, 18'b000000000111001011, 18'b000000000010011010, 18'b111111111110000011, 18'b111111111011100111, 18'b000000000010110000, 18'b000000000000000000, 18'b111111111100001100, 18'b000000000000011011, 18'b000000000001000111, 18'b111111111110100101, 18'b000000000100100010, 18'b111111110000010100, 18'b000000000000101001, 18'b000000000011110100, 18'b111111111111010101, 18'b000000000000001111, 18'b111111111100010001, 18'b111111111111111111, 18'b111111111100110010, 18'b111111111111100111}, 
{18'b000000000011011001, 18'b000000000101100001, 18'b000000001000110011, 18'b111111111100101110, 18'b000000000110101010, 18'b000000000100111001, 18'b000000000000000000, 18'b000000000111010010, 18'b000000000101101101, 18'b111111111110010010, 18'b000000001011001110, 18'b111111111010011010, 18'b000000001001111100, 18'b000000000111001001, 18'b111111101110110101, 18'b111111111111111111, 18'b000000000000000000, 18'b000000000000000101, 18'b000000000100001010, 18'b111111110111111100, 18'b000000000011100010, 18'b111111111100100110, 18'b111111111000001001, 18'b111111111101011111, 18'b000000000101010001, 18'b111111110101011100, 18'b111111111010101110, 18'b111111111111010101, 18'b111111111111111111, 18'b111111110110111110, 18'b000000000110010100, 18'b000000000000000000}, 
{18'b111111111111001101, 18'b000000000000000000, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111010011000, 18'b000000000000001001, 18'b000000000000001000, 18'b111111111111110000, 18'b111111111111100111, 18'b111111111111010000, 18'b000000000010001110, 18'b111111111111111111, 18'b000000000001010100, 18'b111111111010100001, 18'b000000000001101101, 18'b111111111111111111, 18'b000000000010010000, 18'b000000000111001010, 18'b111111111010010110, 18'b000000000000110101, 18'b111111111110011010, 18'b000000000010000011, 18'b000000000011000010, 18'b111111111110101000, 18'b111111111011111110, 18'b000000000000010101, 18'b000000001101010001, 18'b111111111111100111, 18'b111111111111110000, 18'b000000000101001100, 18'b000000000000000000, 18'b000000001101110010}, 
{18'b111111110111101001, 18'b000000000000100101, 18'b111111111100100010, 18'b000000000110001000, 18'b000000000001110000, 18'b111111111111011111, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111011001001, 18'b111111111111011110, 18'b000000000000000000, 18'b111111110111000111, 18'b000000000000001100, 18'b111111111111010111, 18'b111111111111111101, 18'b111111111111111111, 18'b111111111110001000, 18'b000000000000000101, 18'b000000000000000011, 18'b000000000010100010, 18'b000000000000010001, 18'b000000000000000000, 18'b000000000000000000, 18'b111111111111110111, 18'b000000000000000000, 18'b000000000000010010, 18'b000000001001010011, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111111010110, 18'b000000000010110011, 18'b111111111111100101}, 
{18'b111111111111111110, 18'b111111111101100101, 18'b000000000011010001, 18'b000000000000101000, 18'b111111111010000011, 18'b000000000000000000, 18'b000000000100100100, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111110011011, 18'b000000000001110101, 18'b000000000000010011, 18'b000000000101001011, 18'b111111110111001110, 18'b111111111110011111, 18'b111111111111101110, 18'b000000000011011101, 18'b111111111001110110, 18'b000000000000010101, 18'b111111110011111011, 18'b111111111111101100, 18'b111111111110000110, 18'b111111111111010110, 18'b000000000100101110, 18'b111111111110110011, 18'b111111111011100000, 18'b000000000001011100, 18'b000000000000000000, 18'b000000000110010101, 18'b000000001000010111, 18'b111111111010110000, 18'b111111111000110100}, 
{18'b000000000001000101, 18'b000000000000011010, 18'b111111111001010111, 18'b111111111111000101, 18'b111111111111111111, 18'b000000000000000010, 18'b000000000001101100, 18'b000000000110100101, 18'b000000000000000000, 18'b000000000000010100, 18'b000000000001000111, 18'b111111110111010111, 18'b111111111110111011, 18'b111111110110010101, 18'b000000000111101100, 18'b000000000000000000, 18'b111111111111111111, 18'b111111110101101111, 18'b111111111111111111, 18'b111111111110110011, 18'b111111111111101010, 18'b000000000000000000, 18'b000000000000111111, 18'b111111111101100110, 18'b000000000000110110, 18'b000000000110100100, 18'b000000000110110100, 18'b000000000110001111, 18'b000000000100111011, 18'b000000000000000000, 18'b000000000001110100, 18'b000000001100100010}, 
{18'b111111111111100110, 18'b111111111100001100, 18'b000000000110001110, 18'b111111111110010110, 18'b000000000001000111, 18'b000000000010101011, 18'b111111111111111111, 18'b111111111011011010, 18'b111111111110101000, 18'b111111110110011000, 18'b000000000111001010, 18'b000000000000000011, 18'b000000000110101101, 18'b000000001010101110, 18'b111111111110001000, 18'b111111110010000100, 18'b111111111110010101, 18'b000000000111100001, 18'b111111111011011110, 18'b111111111100101010, 18'b000000000000111100, 18'b000000000000000001, 18'b111111110111010001, 18'b111111111100111100, 18'b111111111111010111, 18'b111111111110000011, 18'b000000000001110010, 18'b000000001011010000, 18'b000000000011111011, 18'b111111111111111111, 18'b000000000001010010, 18'b000000000000011100}, 
{18'b000000000000101011, 18'b000000000111010000, 18'b000000000000000000, 18'b000000000100101110, 18'b000000001101010011, 18'b111111111101010001, 18'b111111111111111111, 18'b111111111111010010, 18'b000000000100101100, 18'b111111111100111011, 18'b111111111111111110, 18'b000000000101010101, 18'b000000000000001000, 18'b000000000000011100, 18'b111111100111100100, 18'b111111111110101110, 18'b000000000000000000, 18'b000000000011001101, 18'b111111111111111100, 18'b000000000100110001, 18'b111111111111111111, 18'b111111111101001111, 18'b111111110111000000, 18'b000000000010000101, 18'b000000000100100100, 18'b111111101110010000, 18'b111111111111111111, 18'b000000000000000000, 18'b000000001000101101, 18'b111111110011001011, 18'b000000000000000001, 18'b111111111111111001}, 
{18'b000000000000001001, 18'b111111111010100100, 18'b000000000000110111, 18'b111111111111110000, 18'b000000000000110101, 18'b000000001000011101, 18'b111111110100011001, 18'b000000000000100011, 18'b000000000110110001, 18'b111111111010100110, 18'b111111111111101000, 18'b000000000000110010, 18'b111111111111110110, 18'b000000000010110111, 18'b000000000001101101, 18'b111111111111101110, 18'b000000000001000100, 18'b000000000000000000, 18'b000000000000010110, 18'b000000000110000100, 18'b111111111111100011, 18'b111111111000010000, 18'b111111110110010100, 18'b111111111100111001, 18'b111111110110100011, 18'b000000000011010101, 18'b000000001001111110, 18'b000000000101111001, 18'b111111111111110101, 18'b111111111010000010, 18'b111111111011000001, 18'b000000000000111101}, 
{18'b000000000000110101, 18'b111111111000010110, 18'b111111111111101110, 18'b000000000010011010, 18'b111111111000010110, 18'b000000000010101101, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111111111111, 18'b000000000000000000, 18'b000000000100001110, 18'b111111111111101110, 18'b000000000000001001, 18'b000000000000000000, 18'b000000000010000010, 18'b111111111111101110, 18'b000000000000000010, 18'b111111111111111111, 18'b111111111010110110, 18'b111111110111111010, 18'b111111111111111111, 18'b111111110111011101, 18'b111111111011001011, 18'b111111111010000011, 18'b000000001110001111, 18'b000000000000010010, 18'b111111111111010000, 18'b000000000101000100, 18'b000000001110010111, 18'b000000000110010100, 18'b111111101111000010, 18'b111111111101000010}, 
{18'b000000000110000000, 18'b111111111111111111, 18'b000000000100000001, 18'b111111111111101011, 18'b000000000111101111, 18'b111111111101101101, 18'b000000000001001000, 18'b000000000110101100, 18'b000000000100010010, 18'b111111110111101001, 18'b111111111111000000, 18'b000000000001111101, 18'b000000000001000110, 18'b111111111111110001, 18'b000000000001010110, 18'b000000000000000000, 18'b000000000101110011, 18'b000000000000100011, 18'b000000000101111111, 18'b111111111110111100, 18'b111111111101111101, 18'b111111111110110011, 18'b111111111111111111, 18'b000000000100110101, 18'b111111111100110000, 18'b111111111111111001, 18'b000000000000000000, 18'b000000000000000000, 18'b000000000000000000, 18'b000000000100101011, 18'b111111111010110111, 18'b111111111111101000}, 
{18'b111111111111111111, 18'b111111111111100000, 18'b111111111000100011, 18'b000000000100100011, 18'b000000000011100100, 18'b111111111110001111, 18'b111111111111111111, 18'b111111111100010111, 18'b000000000000000110, 18'b111111111111111111, 18'b111111111011001011, 18'b111111111100000011, 18'b000000000111101010, 18'b000000000000000000, 18'b111111111101111101, 18'b111111111111111111, 18'b000000000011011011, 18'b111111111111111111, 18'b111111111111111111, 18'b111111111100100010, 18'b000000000101000011, 18'b000000000000000000, 18'b000000000010011111, 18'b111111111111100010, 18'b000000000010100000, 18'b000000000000000010, 18'b000000000000000000, 18'b000000000011110110, 18'b111111111100111011, 18'b111111111111010000, 18'b000000000010100100, 18'b111111111110010011}, 
{18'b111111111111101110, 18'b111111111011000100, 18'b000000001001100000, 18'b111111111110111101, 18'b000000000011001001, 18'b111111111011011011, 18'b000000000000000000, 18'b000000000000100011, 18'b111111111000010101, 18'b111111111111110010, 18'b111111111110000001, 18'b000000000000111011, 18'b111111111010110000, 18'b000000000010001101, 18'b000000000011001111, 18'b000000000001110000, 18'b000000000001010111, 18'b111111111111011001, 18'b111111110100101010, 18'b111111111111110010, 18'b111111111111000101, 18'b000000000010001111, 18'b111111111110001110, 18'b111111111111111111, 18'b000000000011001010, 18'b111111111111010001, 18'b111111111111110001, 18'b000000000110001110, 18'b111111111001101000, 18'b111111111011010001, 18'b000000000101100111, 18'b000000000000100100}, 
{18'b000000000110111001, 18'b000000000011001110, 18'b000000000000000000, 18'b111111111101011101, 18'b111111111110101111, 18'b111111111111111111, 18'b000000000000000000, 18'b111111111110111001, 18'b111111111110000000, 18'b111111111110000110, 18'b000000000000000000, 18'b000000000010100010, 18'b000000000000000110, 18'b000000000000110110, 18'b111111111111010010, 18'b000000000000000101, 18'b111111111101100010, 18'b000000000000000000, 18'b111111111111101101, 18'b111111111111111111, 18'b000000000000000010, 18'b000000000000111100, 18'b000000000001100011, 18'b000000000000000000, 18'b000000000000000000, 18'b111111110110001110, 18'b111111111100110011, 18'b000000000000000110, 18'b000000000000010100, 18'b000000000000000001, 18'b111111111101001010, 18'b000000000000010101}, 
{18'b000000000011000000, 18'b111111101111010010, 18'b111111111111111111, 18'b111111111110110010, 18'b111111111100010001, 18'b111111111111110110, 18'b000000000000000000, 18'b000000001000110000, 18'b111111111111010011, 18'b111111111111101001, 18'b000000000001010100, 18'b111111110101011011, 18'b000000000000011000, 18'b111111111000111111, 18'b000000001011100011, 18'b111111111111001010, 18'b111111111100011000, 18'b111111110111001111, 18'b111111111111110101, 18'b111111110100101011, 18'b111111110011000010, 18'b111111111111111111, 18'b000000000000000000, 18'b000000000000000000, 18'b000000000011111001, 18'b111111111111110001, 18'b111111111011001110, 18'b111111111110110101, 18'b111111111111101000, 18'b000000000000000000, 18'b111111111111011111, 18'b111111110100110011}
};

localparam logic signed [17:0] bias [32] = '{
18'b000000000100001110,  // 0.5280959606170654
18'b000000000110101110,  // 0.8414360880851746
18'b000000000011001011,  // 0.397830605506897
18'b000000000011010010,  // 0.4105983078479767
18'b111111100010101111,  // -3.657735586166382
18'b111111111000110100,  // -0.8977976441383362
18'b000000001101101001,  // 1.7051936388015747
18'b111111110101110010,  // -1.2765135765075684
18'b111111111011010101,  // -0.5837795734405518
18'b000000010101100110,  // 2.699671983718872
18'b000000000001101111,  // 0.2170683741569519
18'b000000000111000011,  // 0.8814588785171509
18'b111111101010111011,  // -2.634300947189331
18'b111111110000111110,  // -1.877297282218933
18'b000000001101010011,  // 1.6625694036483765
18'b000000010101111101,  // 2.7459704875946045
18'b111111111100001011,  // -0.47838035225868225
18'b000000001101100101,  // 1.6984987258911133
18'b000000000110110101,  // 0.8548859357833862
18'b000000001000000010,  // 1.0045719146728516
18'b000000001011010110,  // 1.4197649955749512
18'b000000000110101010,  // 0.832463800907135
18'b000000000100010110,  // 0.5434179306030273
18'b000000000111011010,  // 0.9277304410934448
18'b111111111101010000,  // -0.3426123857498169
18'b111111111011100001,  // -0.5587119460105896
18'b111111111011000010,  // -0.6208624839782715
18'b111111110101110000,  // -1.2802538871765137
18'b000000000000011110,  // 0.05940237268805504
18'b111111111001011011,  // -0.8213341236114502
18'b000000000111000001,  // 0.8783953189849854
18'b111111111000011001   // -0.949700653553009
};
endpackage