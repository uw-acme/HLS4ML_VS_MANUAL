//Width: 25
//Int: 9
package dense_2_gen;

localparam logic signed [24:0] weights [64][32] = '{
{25'b0000000000100010011011001, 25'b0000000000000001000010010, 25'b1111111111100111101100011, 25'b1111111111111101010011100, 25'b0000000000100001011011011, 25'b0000000000000000000000001, 25'b1111111111101101100001100, 25'b1111111111111111111111000, 25'b1111111111011100111100101, 25'b0000000000001010001101001, 25'b0000000000000000000000100, 25'b1111111111111111010001100, 25'b1111111111111111111100111, 25'b1111111111100110011001101, 25'b1111111111111001100001001, 25'b1111111111011110011111011, 25'b0000000000000000000000000, 25'b1111111111111110010101101, 25'b1111111111100111100111101, 25'b1111111111101011101110101, 25'b0000000000000000000000110, 25'b0000000000000000000000000, 25'b1111111111111110111110010, 25'b1111111111111111101001101, 25'b0000000000000000000000010, 25'b0000000000001100110111010, 25'b0000000000110001011010111, 25'b0000000000010110011011110, 25'b1111111111111111111100011, 25'b0000000000000110011110110, 25'b1111111111001011100110101, 25'b0000000000000000000010100},
{25'b1111111111110011001011001, 25'b1111111111101100001011011, 25'b1111111111101110010010110, 25'b1111111111111000111001101, 25'b1111111111111111010001111, 25'b0000000000000101100000010, 25'b1111111111100011011010110, 25'b0000000000000000101011001, 25'b0000000000000000100111000, 25'b1111111111110111111101000, 25'b0000000000010011111111000, 25'b1111111111111010011100111, 25'b1111111111111000011101110, 25'b1111111111100100001111100, 25'b0000000000000000111101001, 25'b1111111111111001110111000, 25'b0000000000000001100110001, 25'b1111111111100111000100111, 25'b0000000000010101111111011, 25'b0000000000011101011000110, 25'b1111111111111011111111100, 25'b1111111111111111010001111, 25'b1111111111111111111101110, 25'b0000000000000011000001111, 25'b1111111111110110111000001, 25'b0000000000100011001101011, 25'b0000000000011111101100001, 25'b0000000000000001000110000, 25'b0000000000000011101001110, 25'b1111111111000001101100110, 25'b0000000000000000111100010, 25'b0000000000000000000000000},
{25'b0000000000001001010001101, 25'b1111111111110001010100010, 25'b1111111111101111011010011, 25'b1111111111111010101001101, 25'b1111111111110110000101111, 25'b1111111111110101000101100, 25'b1111111111101000010101100, 25'b0000000000000000100100101, 25'b1111111111101110101110010, 25'b0000000000000001001001010, 25'b0000000000000000010001010, 25'b1111111111110101101011001, 25'b0000000000001011100100100, 25'b1111111111110111101111100, 25'b1111111111111111110100111, 25'b1111111111111011010011011, 25'b0000000000000000101000100, 25'b0000000000001100001110100, 25'b0000000000000111100000010, 25'b0000000000011101011010111, 25'b0000000000000101010000101, 25'b1111111111110101001111010, 25'b0000000000000000000011000, 25'b0000000000000100011110010, 25'b1111111111111101101001110, 25'b0000000000011010110010100, 25'b0000000000010011000110010, 25'b0000000000001100011001100, 25'b1111111111111111111100110, 25'b1111111111101100100010000, 25'b1111111111111110010001001, 25'b0000000000001100101101100},
{25'b0000000000010001101011101, 25'b0000000000000010011101010, 25'b0000000000000110110001111, 25'b1111111111111110110000101, 25'b1111111110111110110101111, 25'b0000000000000000000000000, 25'b0000000000000000000010100, 25'b0000000000011100111101000, 25'b0000000000011111000011010, 25'b1111111111111110010011000, 25'b1111111111111111111111111, 25'b0000000000000000000000111, 25'b0000000000000000000010110, 25'b0000000000000000101000001, 25'b1111111111111101101010010, 25'b0000000000011011011111000, 25'b0000000000000000000001010, 25'b1111111111111100110110110, 25'b1111111111111111111111101, 25'b1111111111101001011101100, 25'b1111111111111000001011000, 25'b0000000000000110010101110, 25'b1111111111110111111000011, 25'b1111111111111111111101010, 25'b0000000000000000011111100, 25'b1111111111111001100000001, 25'b0000000000001001010110010, 25'b1111111111111111111110111, 25'b1111111111111111111111000, 25'b1111111111111111111111110, 25'b1111111111100100011101111, 25'b0000000000100111101110000},
{25'b1111111110101000101001110, 25'b1111111111111100110100110, 25'b1111111111111111011110000, 25'b0000000000000000101011100, 25'b1111111111111100101000110, 25'b0000000000000000110110001, 25'b1111111111111001101101100, 25'b1111111111101100110101110, 25'b0000000000000110111100011, 25'b1111111111111101011010110, 25'b1111111111111110010000100, 25'b1111111111111111111110111, 25'b1111111111111111111110111, 25'b0000000000011010111010011, 25'b0000000000000000000000110, 25'b0000000000101010000111111, 25'b1111111111111111111111011, 25'b0000000000011011111011101, 25'b1111111111001100110011011, 25'b0000000000000000000010100, 25'b1111111111110001101101110, 25'b0000000000010101100101000, 25'b0000000000100001000011010, 25'b0000000000000000000000111, 25'b0000000000000101110011100, 25'b0000000000010100110110101, 25'b0000000000011110100011111, 25'b0000000000000010001110000, 25'b1111111111111111011011011, 25'b1111111111111111111110110, 25'b1111111111111110001111000, 25'b0000000000011100111101011},
{25'b0000000000000111011000101, 25'b1111111111111111111110110, 25'b0000000000010011000110101, 25'b1111111110101100111111111, 25'b1111111101001111101110010, 25'b1111111111010011001001100, 25'b0000000000101101010101111, 25'b1111111110110000010111111, 25'b1111111111111111111101100, 25'b1111111110101001010011001, 25'b1111111110111111110111101, 25'b1111111111010100010110000, 25'b0000000000101101001110110, 25'b1111111111111111111111101, 25'b1111111111111110000110011, 25'b0000000000000000000000011, 25'b1111111111111111111111111, 25'b1111111111111111111100110, 25'b1111111111101111000101000, 25'b1111111111111111111111001, 25'b1111111111000001011000100, 25'b0000000000000000000000001, 25'b0000000000010111110011010, 25'b1111111111111111111111100, 25'b0000000000000010110100011, 25'b0000000000100010010001001, 25'b0000000000000110100011111, 25'b1111111111111111111111111, 25'b1111111111111111111111001, 25'b0000000000011010010100000, 25'b1111111111111011101000011, 25'b0000000000011001101011001},
{25'b1111111111111011011001010, 25'b1111111111101011110111111, 25'b1111111111100001000100100, 25'b1111111111111001111111011, 25'b1111111111011011000100010, 25'b0000000000001000011101111, 25'b1111111111101000111101111, 25'b1111111111101101110100111, 25'b1111111111001010111010010, 25'b0000000000000110001100101, 25'b1111111111111111010110011, 25'b1111111111101011101000000, 25'b0000000000001111001110111, 25'b1111111111111110101101000, 25'b1111111111111010101100010, 25'b1111111110111001001000000, 25'b1111111111111111111110010, 25'b0000000000001010110000001, 25'b0000000000011000100010010, 25'b1111111111101011001110100, 25'b1111111111101100110011101, 25'b1111111111110111111111001, 25'b1111111111111111110101011, 25'b0000000000000011100010010, 25'b1111111111111010001011101, 25'b1111111110101101000010011, 25'b1111111111011110000101110, 25'b1111111111111010001111101, 25'b0000000000000000101110111, 25'b1111111111111101010001100, 25'b0000000000000011111010101, 25'b1111111111111111111010001},
{25'b1111111111101100010110000, 25'b1111111111110100011011010, 25'b1111111111110101110101001, 25'b1111111111100001101000110, 25'b1111111111110001001011011, 25'b1111111111111111111101101, 25'b0000000000001101010111110, 25'b1111111111110101111000010, 25'b0000000000011001101011100, 25'b0000000000000000000001010, 25'b0000000000000000000001000, 25'b1111111111111111111111000, 25'b0000000000011100000001000, 25'b0000000000000000000001001, 25'b1111111111111111111110100, 25'b1111111111110110111100011, 25'b1111111111111111111101000, 25'b0000000000000000000000100, 25'b1111111111111111111100110, 25'b0000000000000000000000111, 25'b1111111111111111111101001, 25'b1111111111111111111011110, 25'b0000000000000000000001101, 25'b1111111111111111111111111, 25'b0000000000000101101001100, 25'b1111111111101000111101110, 25'b0000000000000001110001100, 25'b1111111111111111111110000, 25'b1111111111110110110001100, 25'b1111111111111111111010011, 25'b0000000000000000000011110, 25'b1111111111111111111110110},
{25'b1111111111000010111000110, 25'b1111111111111000101100000, 25'b1111111111001111010110010, 25'b0000000000001111101001111, 25'b0000000000111110010101001, 25'b1111111111111111111111111, 25'b1111111111111100010010010, 25'b0000000000011110100101010, 25'b1111111111000111110101100, 25'b1111111111111010000001100, 25'b0000000000000000000001000, 25'b1111111111100110001101100, 25'b1111111111111111111101001, 25'b0000000000001001101111111, 25'b1111111111100111100111100, 25'b0000000001100000100000000, 25'b1111111111111110111001111, 25'b0000000000000101111111010, 25'b0000000000011010100101111, 25'b0000000000011111010110000, 25'b0000000000000000000001110, 25'b1111111111010101000001000, 25'b0000000000000000000001110, 25'b0000000000110100101011101, 25'b1111111111101000110011111, 25'b0000000001011001010011001, 25'b1111111111101100111001100, 25'b1111111111100101111001111, 25'b1111111111000011100101111, 25'b1111111111000100100101100, 25'b0000000000000000000010100, 25'b0000000000000110110101110},
{25'b0000000000000000000001000, 25'b1111111111111110000001001, 25'b1111111111110110100011000, 25'b0000000000000000000000010, 25'b0000000000100111011111100, 25'b1111111111111101011010110, 25'b1111111111110111110110110, 25'b0000000000001011110000011, 25'b0000000000001100111111001, 25'b0000000000000000011100001, 25'b1111111111111110111010001, 25'b1111111111111111111101001, 25'b1111111111111111111111111, 25'b1111111111110001011101010, 25'b1111111111111111111111010, 25'b0000000000000000000010001, 25'b0000000000000000000000001, 25'b1111111111111111010110110, 25'b0000000000000000010001101, 25'b0000000000001010110111110, 25'b0000000000000010011101110, 25'b1111111111111111111111010, 25'b0000000000000000000001111, 25'b0000000000000000111010110, 25'b0000000000000100111010010, 25'b1111111111101111000110100, 25'b0000000000001000101100111, 25'b0000000000011111110100011, 25'b1111111111111111111111110, 25'b0000000000000000110010000, 25'b0000000000000110010110001, 25'b0000000000001000111000111},
{25'b0000000000001100010100101, 25'b0000000000000000000000011, 25'b1111111111110010110011100, 25'b1111111111011111111001010, 25'b1111111110011010010111001, 25'b0000000000010001000010000, 25'b0000000000000000000011101, 25'b1111111110010110000110001, 25'b0000000000000100101001111, 25'b1111111111111111111101101, 25'b0000000000000000011110001, 25'b1111111111111111110010101, 25'b0000000000000001010110100, 25'b0000000000000000000010000, 25'b1111111111111101100101001, 25'b1111111111001111001001100, 25'b1111111111111111111111000, 25'b0000000000011100001001010, 25'b0000000000010000001011011, 25'b0000000000011000011110110, 25'b1111111111000111101110101, 25'b1111111111010010011100110, 25'b0000000000001111010111101, 25'b1111111111111011100010101, 25'b1111111111111010000110011, 25'b0000000000101101111001000, 25'b1111111111110011101000011, 25'b1111111111111111111101110, 25'b1111111111111111111110111, 25'b0000000000011011000001100, 25'b1111111111111111111110110, 25'b0000000000000000110011100},
{25'b1111111111100110101111101, 25'b1111111111000000111001010, 25'b0000000000000000000000000, 25'b1111111111111111101110101, 25'b0000000000101010100000011, 25'b1111111111011101100011000, 25'b1111111111100011101010011, 25'b0000000000001110110101101, 25'b1111111111111111111011001, 25'b0000000000010011000010101, 25'b0000000000001001011110100, 25'b1111111111110110010100010, 25'b0000000000000000000010001, 25'b0000000000000001110011111, 25'b1111111111111101010010011, 25'b1111111111011111100111010, 25'b0000000000010110011101001, 25'b0000000000000011101001110, 25'b0000000000100110000011001, 25'b0000000000001011000101000, 25'b0000000000000000000000100, 25'b1111111111111011001010010, 25'b0000000000010000001000100, 25'b1111111111110100111100001, 25'b1111111111011000100100101, 25'b1111111111111111001001001, 25'b0000000000010111101011110, 25'b1111111111111111111110010, 25'b0000000000000001000101000, 25'b1111111111110011111000010, 25'b0000000000010001100110100, 25'b0000000000100011010111001},
{25'b0000000000000001111100001, 25'b0000000000000000000001000, 25'b0000000000011100000100100, 25'b0000000000000001000100111, 25'b1111111111111010110010101, 25'b0000000000010111000110011, 25'b0000000000001011110011101, 25'b1111111111111111111101100, 25'b0000000000000000000110101, 25'b1111111111101110000011100, 25'b1111111111111001000000010, 25'b1111111111101010100101000, 25'b1111111111111111111110001, 25'b0000000000000110011101010, 25'b1111111111110111001011011, 25'b0000000001101011111011010, 25'b0000000000000000000010010, 25'b1111111111110011111101001, 25'b1111111111100111110110011, 25'b1111111111111110010100000, 25'b0000000000011001011011101, 25'b0000000000010000011000010, 25'b0000000000000000000001101, 25'b1111111111111111101011010, 25'b0000000000011100000110100, 25'b0000000000100010010100101, 25'b0000000000111111011001110, 25'b0000000000000001010100111, 25'b0000000000000000000001010, 25'b0000000000000000000011101, 25'b1111111111111110011110011, 25'b1111111111110110110110001},
{25'b1111111111101100000000111, 25'b0000000000000110001100011, 25'b0000000000000101000010101, 25'b1111111111100000010110111, 25'b1111111111011101100000000, 25'b0000000000111100000001101, 25'b0000000000000110010010101, 25'b0000000000000000000000001, 25'b1111111111101011011011001, 25'b1111111111110100101100110, 25'b0000000000010000100101000, 25'b0000000000001001000100011, 25'b0000000000000000000100101, 25'b1111111111110101111101100, 25'b0000000000100100100111100, 25'b1111111111111111111110010, 25'b1111111111111110010000110, 25'b0000000000000000000001010, 25'b0000000000000001101011100, 25'b1111111111111010000011001, 25'b0000000000001010000001100, 25'b0000000000000010000001001, 25'b0000000000001110100110101, 25'b1111111111111111111110000, 25'b0000000000000000011011100, 25'b0000000001010100001111001, 25'b1111111111111000110010001, 25'b1111111111111101000011101, 25'b1111111111111111111110111, 25'b1111111111110010000001001, 25'b1111111111111010110111110, 25'b0000000000010110100001100},
{25'b0000000000000111100010110, 25'b0000000000001001011111101, 25'b0000000000101001110010100, 25'b1111111111111010111010011, 25'b0000000000001100111011001, 25'b0000000000101100111010010, 25'b0000000000000000000101100, 25'b1111111111111100001111010, 25'b0000000000001111000110101, 25'b1111111111110001011011100, 25'b1111111111111111111111001, 25'b1111111111110000101111111, 25'b0000000000000000000010101, 25'b0000000000110010010101000, 25'b1111111111111101101111011, 25'b0000000000000000001101001, 25'b0000000000011110001110110, 25'b0000000000000000000101100, 25'b0000000000000000011000010, 25'b1111111111010111111101010, 25'b1111111111100000100100101, 25'b1111111111111011011000100, 25'b1111111111111111111111110, 25'b1111111111101101010100111, 25'b1111111111111011011000011, 25'b1111111111110101011100110, 25'b1111111111100110110111000, 25'b1111111111100100110011110, 25'b0000000000000011110110001, 25'b0000000000001110010010011, 25'b1111111111001101001001110, 25'b0000000000000000011010100},
{25'b1111111111011001110010111, 25'b0000000000000000000000111, 25'b1111111111111110000110011, 25'b1111111111111001101001010, 25'b1111111111111111111110000, 25'b0000000000010001000100010, 25'b1111111111110110000110001, 25'b0000000000100010101100010, 25'b1111111111010001100001001, 25'b1111111111111111111011010, 25'b0000000000000000000000011, 25'b1111111111111111111111111, 25'b0000000000000000000011000, 25'b0000000000000000000001001, 25'b1111111111111111100010000, 25'b1111111111110100011001111, 25'b0000000000001010001001000, 25'b0000000000010111011101010, 25'b1111111111111110110100000, 25'b1111111111011111110101110, 25'b1111111111111000011110101, 25'b0000000000001110010100001, 25'b0000000000001000000100000, 25'b0000000000000000000011111, 25'b0000000000000000011001000, 25'b0000000000001010011101001, 25'b1111111111100001010110100, 25'b0000000000000000000000111, 25'b1111111111111111111111101, 25'b0000000000000000011011000, 25'b0000000000000000000100001, 25'b1111111111101111111001101},
{25'b1111111111010100111110011, 25'b1111111111111111010000010, 25'b1111111111111111100111101, 25'b1111111111111101110001101, 25'b1111111111111111011000100, 25'b0000000000001101100000010, 25'b0000000000000000110110010, 25'b0000000000000100011100000, 25'b0000000000000100111000101, 25'b0000000000001000000011101, 25'b0000000000001010000110010, 25'b0000000000010100101000011, 25'b0000000000000011011011100, 25'b1111111111110011100111110, 25'b0000000000000000000100000, 25'b0000000000110000110101000, 25'b0000000000000000000010101, 25'b0000000000000000001001001, 25'b1111111111111111101011010, 25'b0000000000001110000101100, 25'b0000000000010010001110010, 25'b0000000000000011111100111, 25'b0000000000000101010001101, 25'b1111111111111100001100110, 25'b1111111111111011111000100, 25'b0000000000000011011001011, 25'b1111111111110111011010101, 25'b1111111111101111110010100, 25'b0000000000011010110100001, 25'b1111111111111100000100001, 25'b0000000000000100000011011, 25'b1111111111100111111101101},
{25'b0000000000000000000001001, 25'b1111111111111111111111110, 25'b0000000000000100110100101, 25'b0000000000000000000001001, 25'b0000000001110100000011110, 25'b1111111111111111111010000, 25'b0000000000000000000000001, 25'b1111111111111111111111111, 25'b0000000000001110000010010, 25'b1111111111110110011000101, 25'b0000000000000000000000001, 25'b0000000000000000000000101, 25'b0000000000000000001001001, 25'b0000000000010000100001110, 25'b0000000000000000000000011, 25'b1111111111101101011001010, 25'b1111111111111111111111011, 25'b1111111111110111011011010, 25'b0000000000101001111010011, 25'b0000000000000000000001111, 25'b1111111111111111111111111, 25'b1111111111111111111101101, 25'b0000000000000000000000110, 25'b1111111111111111111111111, 25'b0000000000000000000000010, 25'b0000000000001000101111111, 25'b0000000000000000000000011, 25'b0000000000000000000000100, 25'b1111111111111111111111111, 25'b1111111111111111111110111, 25'b0000000000000000000001111, 25'b0000000000000101010011010},
{25'b1111111111111111100100100, 25'b0000000000000011101101110, 25'b1111111111111111111001111, 25'b0000000000000110001000011, 25'b1111111111111010010100001, 25'b1111111111110000101110110, 25'b1111111111111000000000111, 25'b0000000000100011100011111, 25'b0000000000000000000010011, 25'b0000000000001100011001100, 25'b1111111111111110100101101, 25'b0000000000001000010011111, 25'b1111111111111011110000010, 25'b1111111111101011110101011, 25'b1111111111100111100111010, 25'b0000000000000001101011010, 25'b1111111111111111111111111, 25'b1111111111111011100010101, 25'b0000000000000000000000110, 25'b0000000000000000000011100, 25'b1111111111111111111011110, 25'b0000000000001001101100011, 25'b0000000000000100100100000, 25'b1111111111101111111001100, 25'b0000000000001110010011100, 25'b1111111111101010111100101, 25'b0000000000000000010001111, 25'b0000000000000000000000000, 25'b1111111111101010100010101, 25'b0000000000000000000000011, 25'b0000000000000101110101101, 25'b1111111111111100000001100},
{25'b1111111111111110100001110, 25'b1111111111110011010101011, 25'b0000000000000000000001111, 25'b1111111111111000010110010, 25'b0000000000011011101001001, 25'b1111111111111111111101101, 25'b1111111111111101010101001, 25'b0000000000001101101010100, 25'b1111111111001101111110100, 25'b0000000000000000000001000, 25'b1111111111111011000100001, 25'b1111111111111111101110101, 25'b0000000000101100111111100, 25'b0000000000011101010111100, 25'b1111111111110011010010110, 25'b1111111111111101010101111, 25'b1111111111111111111101111, 25'b0000000000000000000101100, 25'b1111111111111111111110101, 25'b0000000000000000000010110, 25'b0000000000000000000001100, 25'b1111111111101110100111111, 25'b1111111111110000110001101, 25'b0000000000010000110000001, 25'b0000000000000000000000011, 25'b1111111111101110011101010, 25'b0000000000000011001000010, 25'b1111111111110101101101111, 25'b1111111111111011101111100, 25'b0000000000010001011001100, 25'b0000000000000000000100101, 25'b1111111111100000010111111},
{25'b0000000001010001001111110, 25'b0000000000101011110001011, 25'b1111111111100000000101101, 25'b0000000000000000011010101, 25'b1111111111010011101101010, 25'b0000000000000000000000100, 25'b0000000000011100100001011, 25'b0000000000000011111110110, 25'b0000000000011100101001011, 25'b1111111111111111111101101, 25'b1111111111101100001011110, 25'b1111111111110101111101000, 25'b0000000000010010001001010, 25'b0000000000000011100010110, 25'b1111111111110011011011110, 25'b0000000000010000110111001, 25'b0000000001000100100000110, 25'b1111111111101111010111000, 25'b1111111111011010000110100, 25'b0000000000000000000000110, 25'b1111111111111100010101001, 25'b1111111111101001011001001, 25'b1111111111111110011100111, 25'b1111111111111111110011100, 25'b0000000000001011000000010, 25'b1111111111010001110111100, 25'b0000000000001011011000100, 25'b1111111111111111110111001, 25'b0000000000000000000010101, 25'b0000000000001101111101011, 25'b1111111111111100010011110, 25'b0000000000000111101000000},
{25'b1111111111110100001001111, 25'b1111111111100111011011111, 25'b1111111111111011010110111, 25'b1111111111101010100101011, 25'b1111111111111101110011100, 25'b0000000000000110010011010, 25'b0000000000000000000001110, 25'b1111111111111110100011000, 25'b0000000000000100110100011, 25'b1111111111111111100011110, 25'b0000000000000000000001111, 25'b1111111111100100001110111, 25'b0000000000001101000011101, 25'b0000000000001010010010100, 25'b1111111111110010111001101, 25'b0000000000111000110001000, 25'b1111111111111111111110001, 25'b0000000000000000000001101, 25'b1111111111111111011111000, 25'b0000000000000000000000101, 25'b0000000000101000011101001, 25'b1111111111000011110000111, 25'b1111111111110010001000111, 25'b1111111111111000110101110, 25'b1111111111111101100111101, 25'b0000000000011001001110110, 25'b1111111111111001010010110, 25'b0000000000000010010000011, 25'b0000000000111101111111100, 25'b1111111110111110011001100, 25'b1111111111010001000000100, 25'b0000000000000010110111111},
{25'b0000000000000010001001110, 25'b1111111111111000011110001, 25'b1111111111111111111111111, 25'b0000000000000000000001110, 25'b1111111110100011111110110, 25'b1111111110110010011000100, 25'b0000000000000000001100011, 25'b1111111111111111111110111, 25'b1111111111011110000100101, 25'b0000000000000011001010000, 25'b0000000000000000000000011, 25'b1111111111111100011110110, 25'b0000000000000000000000001, 25'b1111111111111000100010000, 25'b1111111111111001010001000, 25'b1111111111110111001100000, 25'b1111111111101101001011111, 25'b0000000000100100001000011, 25'b0000000000000000000000111, 25'b0000000000000101111010011, 25'b1111111111111111111100100, 25'b1111111111110110111110001, 25'b0000000000000000000000101, 25'b1111111111110100111001001, 25'b0000000000011100000110100, 25'b1111111110110000010101010, 25'b0000000000011100001011001, 25'b1111111111111111111111000, 25'b1111111111111111011000011, 25'b0000000000011001100110111, 25'b1111111111111111111111010, 25'b0000000000011110001111101},
{25'b1111111111111111111110100, 25'b0000000000000000101010011, 25'b1111111111111010011110101, 25'b0000000000001001100111100, 25'b0000000000000111000101100, 25'b1111111111010100001110111, 25'b0000000000000000000010000, 25'b0000000000001000001111101, 25'b0000000001001010001100010, 25'b1111111111111110110110101, 25'b0000000000000000000000001, 25'b0000000000000111001101101, 25'b0000000000101101111100110, 25'b1111111111111011111100000, 25'b0000000000000001110010100, 25'b0000000000001100111011100, 25'b1111111111111111111111001, 25'b0000000000000011100011100, 25'b1111111111111111111101110, 25'b0000000000000000000111101, 25'b1111111111011100111101110, 25'b0000000000000100111010001, 25'b0000000000001000111111101, 25'b0000000000000010111010001, 25'b1111111111111111111110111, 25'b0000000000011011111100001, 25'b0000000000000000100100111, 25'b0000000000010000001000101, 25'b1111111111001010100011001, 25'b0000000000001101001010010, 25'b0000000000110010101001100, 25'b0000000000000000101110010},
{25'b1111111111010011000101010, 25'b0000000000011011000001001, 25'b1111111111011110101010100, 25'b0000000000001111101111010, 25'b1111111111110010100000011, 25'b0000000000000000000010001, 25'b0000000000111111101100111, 25'b1111111111100010001101010, 25'b1111111111011010101110101, 25'b0000000000010101111011110, 25'b1111111111100011011111111, 25'b1111111111111100111111010, 25'b1111111111111111111001000, 25'b0000000000101100000010011, 25'b1111111111111111110011010, 25'b1111111111011001011000010, 25'b1111111111111111111111011, 25'b0000000000111000011011110, 25'b1111111111000011101101110, 25'b1111111111111100111001010, 25'b0000000000101000100001111, 25'b1111111111010001100101000, 25'b0000000000000110110010001, 25'b1111111111111110000100010, 25'b0000000000100010101111101, 25'b1111111110111110111001011, 25'b1111111111010001100100010, 25'b1111111111100110111001010, 25'b1111111111111111111111011, 25'b0000000000001101010000001, 25'b0000000000000011001101110, 25'b0000000000010110110101001},
{25'b1111111111110100011000110, 25'b0000000000000110101010000, 25'b1111111111111111111110110, 25'b0000000000010011001011010, 25'b1111111111111011001001011, 25'b0000000000011101000011101, 25'b0000000000000000010000010, 25'b1111111111111110100100011, 25'b1111111111111111101111001, 25'b0000000000000000001001011, 25'b0000000000000000000000101, 25'b1111111111111111111111111, 25'b1111111111111111110001000, 25'b0000000001000010100101010, 25'b0000000000000001100111010, 25'b0000000000011000001011000, 25'b0000000000000000000010010, 25'b1111111111100100111010011, 25'b1111111111110110001110110, 25'b1111111111111111111111011, 25'b1111111111111101111000010, 25'b0000000000000101011001001, 25'b1111111111111111111111011, 25'b1111111111101000010011000, 25'b1111111111111111111111011, 25'b0000000000100101110101101, 25'b0000000000100111101101100, 25'b1111111111111111111111101, 25'b1111111111111101111010100, 25'b0000000000000000000000010, 25'b1111111111111111111011111, 25'b1111111111110011101010000},
{25'b1111111111110101101010100, 25'b0000000000000000000000110, 25'b0000000000100010111100001, 25'b0000000000000000000000101, 25'b0000000000000000000001000, 25'b1111111111110001011101111, 25'b0000000000000000000011000, 25'b1111111110010001011100000, 25'b0000000000011011100101101, 25'b0000000000000001110000100, 25'b0000000000000011011010111, 25'b1111111111010001111100000, 25'b0000000000000000011100000, 25'b1111111111101110011010011, 25'b1111111111111011110000001, 25'b0000000000000000000001011, 25'b0000000000000010100000111, 25'b0000000000000000000001101, 25'b0000000000001110011000110, 25'b0000000000000000000010010, 25'b1111111111111110110111010, 25'b0000000000101010001001000, 25'b0000000000110000001100011, 25'b1111111111100011101110010, 25'b1111111111101101110100100, 25'b0000000000011111111100011, 25'b1111111111011000111000010, 25'b0000000000000011110000100, 25'b1111111111111111111011001, 25'b1111111111111111111111001, 25'b1111111111111111111110011, 25'b0000000000010111100100110},
{25'b1111111111110001011110010, 25'b1111111111111111111011100, 25'b1111111111100001011000100, 25'b1111111111100110001001010, 25'b1111111111111110001111010, 25'b1111111111101110101111010, 25'b0000000000000000000000101, 25'b0000000000001011101010001, 25'b1111111111100001010100101, 25'b1111111111110101010101110, 25'b1111111111111001101001101, 25'b0000000000000000000010000, 25'b0000000000000011100100111, 25'b1111111111111110101111011, 25'b1111111111111000001100100, 25'b0000000000001100001111010, 25'b0000000000011100100001111, 25'b0000000000010000110010110, 25'b1111111111101111010000111, 25'b0000000000000110001111101, 25'b1111111111111110011111110, 25'b1111111111111100010110010, 25'b0000000000000010111000100, 25'b0000000000000010000010010, 25'b1111111111110111000111010, 25'b0000000000001011011001111, 25'b1111111111110100011001010, 25'b0000000000000111101010000, 25'b1111111111111111111110001, 25'b1111111111011010001101010, 25'b1111111111111100101000100, 25'b0000000000011100110010011},
{25'b1111111111111100100011101, 25'b1111111111110101011010010, 25'b0000000000001001110110011, 25'b0000000000100000011001110, 25'b0000000000001010110110100, 25'b0000000000001010100011000, 25'b0000000000000101111110100, 25'b1111111111100110001110000, 25'b1111111111100101101111000, 25'b0000000000001000110001000, 25'b0000000000000001100011011, 25'b0000000000000101100001111, 25'b0000000000000010110111000, 25'b0000000000000000101100100, 25'b0000000000011010010000110, 25'b0000000000000000111100001, 25'b1111111111111001000110011, 25'b0000000000001101001110101, 25'b1111111111111100001101010, 25'b1111111111111011011011011, 25'b0000000000001110000101111, 25'b1111111111110000001000111, 25'b1111111111111100100101110, 25'b0000000000010000010000011, 25'b0000000000000010110101110, 25'b1111111111110010010110001, 25'b1111111111100110101011010, 25'b1111111111111110011111110, 25'b1111111111011100010001010, 25'b0000000000000111101100001, 25'b0000000000001101000001001, 25'b0000000000000000001001111},
{25'b1111111111111110010000101, 25'b1111111111111101011110011, 25'b1111111111111110011110111, 25'b1111111111111011100100001, 25'b1111111111101111001010011, 25'b1111111111101110000010111, 25'b0000000000001000000101011, 25'b0000000000000001000011110, 25'b1111111111101000101001010, 25'b0000000000010101011011010, 25'b1111111111111101010101101, 25'b1111111111111111111011010, 25'b1111111111110001111001110, 25'b0000000000000000101010111, 25'b0000000000000011110001111, 25'b1111111111111001010001000, 25'b1111111111111101111101111, 25'b1111111111111010101010011, 25'b1111111111110101101101110, 25'b0000000000000000000010011, 25'b1111111111101110000001111, 25'b0000000000001101000010111, 25'b1111111111100100111011110, 25'b0000000000000000101001000, 25'b0000000000000101010111111, 25'b0000000000001111110111100, 25'b0000000000000011011001111, 25'b0000000000000000110001001, 25'b0000000000100101011000000, 25'b0000000000000110100110110, 25'b0000000000000000000010010, 25'b0000000000001010101110110},
{25'b1111111111111101100001011, 25'b0000000000100000010110100, 25'b1111111111111111111111010, 25'b1111111111111011110010010, 25'b1111111111100100101001011, 25'b1111111111110110011000110, 25'b0000000000110100101010100, 25'b1111111110100111110010111, 25'b1111111111010011010000001, 25'b1111111111100110011101100, 25'b1111111111100011111010010, 25'b1111111111011111100011001, 25'b1111111111111111111011011, 25'b0000000000111101111111100, 25'b1111111111111100101001110, 25'b0000000000000000000001000, 25'b1111111111100100111110000, 25'b0000000000111001000011011, 25'b1111111111001011001010101, 25'b0000000000000000000001010, 25'b1111111111111111111101101, 25'b1111111111010100111101111, 25'b0000000000000000000001011, 25'b1111111111111111111111111, 25'b0000000000000111001100011, 25'b1111111111111000101010000, 25'b1111111111101101000101110, 25'b1111111111111111111111110, 25'b0000000000010110010110000, 25'b0000000000000000011011111, 25'b1111111111110101101110110, 25'b0000000000000000000110111},
{25'b0000000000101111000110100, 25'b1111111111110001101011111, 25'b0000000000010000111000110, 25'b1111111111111011110111011, 25'b0000000000001001110001000, 25'b1111111111111111100001111, 25'b1111111111111111101000100, 25'b1111111111110100000110110, 25'b0000000000000000000010011, 25'b0000000000001011110011001, 25'b1111111111111111111111111, 25'b1111111111111000011111001, 25'b1111111111111111111100011, 25'b0000000000011101010001000, 25'b0000000000000010011101110, 25'b0000000000000101001011010, 25'b0000000000000011000100001, 25'b1111111111111100111011100, 25'b0000000000000010100110001, 25'b0000000000000000000001100, 25'b1111111111111110110110001, 25'b1111111111111111111111101, 25'b1111111111011000111000001, 25'b1111111111111111111111010, 25'b0000000000000111011001111, 25'b1111111111110001000111110, 25'b1111111111101110101100110, 25'b1111111111111111111111100, 25'b1111111111111111111001011, 25'b0000000001000111011001010, 25'b1111111111011011011011101, 25'b1111111111110001001000110},
{25'b1111111111111010010111010, 25'b1111111111110010110010001, 25'b1111111111110111101111111, 25'b0000000000000100101001010, 25'b0000000000010001110111000, 25'b1111111111101111011000011, 25'b1111111111111111110101011, 25'b1111111111100011110111000, 25'b0000000000000111110001101, 25'b0000000000010001011010010, 25'b1111111111100100101100000, 25'b1111111111011111101001010, 25'b0000000000000011000011100, 25'b1111111110101000100001110, 25'b1111111111110110010110110, 25'b1111111111110000001100011, 25'b1111111111100110101011110, 25'b1111111111111111111101010, 25'b0000000000010001001011110, 25'b0000000000000000000000011, 25'b1111111111111010001010001, 25'b1111111111111010010010110, 25'b0000000000000000000000011, 25'b0000000000000000000000111, 25'b1111111111111000011100111, 25'b1111111110011111011100101, 25'b1111111110111000111010110, 25'b1111111111011101000111101, 25'b0000000000000111001010010, 25'b0000000000011010011001111, 25'b1111111111111111111110000, 25'b0000000000011110110000110},
{25'b1111111111110100001101010, 25'b1111111111100100100000001, 25'b0000000000010100111101011, 25'b0000000000001001100011001, 25'b0000000000000101100011110, 25'b1111111111110100001111000, 25'b1111111111111011110100110, 25'b0000000000001100100111110, 25'b0000000001000100111111111, 25'b1111111111101010000101100, 25'b1111111111111111111111100, 25'b1111111111111111111111101, 25'b0000000000001111000011100, 25'b1111111111111000111110010, 25'b1111111111111101101101110, 25'b1111111111111101110111011, 25'b1111111111110011001101110, 25'b1111111111111111111001000, 25'b0000000000000000000000011, 25'b0000000000011101000000101, 25'b1111111111101110111111000, 25'b1111111111111111100111110, 25'b0000000000010000011101110, 25'b1111111111111110101100110, 25'b0000000000000000000000101, 25'b0000000001000011010111110, 25'b0000000000101001100000001, 25'b0000000000000000011010011, 25'b0000000000000000000010111, 25'b1111111111001010001000101, 25'b1111111111110111010000101, 25'b1111111111111111111111111},
{25'b0000000000000001111011011, 25'b0000000000000110001100000, 25'b1111111111111110001111011, 25'b0000000000000000000000101, 25'b0000000000011101100111111, 25'b1111111111000010001001111, 25'b0000000000000000000001010, 25'b1111111111110011110101100, 25'b0000000000010111110111100, 25'b0000000000000000000000110, 25'b1111111111111101101000100, 25'b0000000000000000000000111, 25'b0000000000000000000010110, 25'b1111111111111111111110100, 25'b0000000000000000101111110, 25'b1111111111110010001111110, 25'b0000000000100001001101111, 25'b1111111111111111010011001, 25'b1111111111111110000001110, 25'b1111111111111111111111111, 25'b0000000000000000000010110, 25'b1111111111111111000010000, 25'b0000000000000000000010001, 25'b1111111111111111111111101, 25'b0000000000000001101001011, 25'b1111111111010111011011101, 25'b0000000000000110100111011, 25'b0000000000010111011101000, 25'b1111111111111111100101111, 25'b0000000000001100000100000, 25'b1111111111111111111101011, 25'b0000000000001001100100111},
{25'b1111111111100110001111111, 25'b0000000000000001001010111, 25'b1111111111000010010000100, 25'b0000000000000000111000101, 25'b1111111111111001100110111, 25'b1111111111111010111010010, 25'b1111111111111111110110000, 25'b1111111111110100010101110, 25'b1111111111111011011001100, 25'b1111111111110111101000111, 25'b0000000000000110000001010, 25'b0000000000000011011100010, 25'b1111111111101001010011101, 25'b0000000000000000000100011, 25'b1111111111111111110000111, 25'b1111111111111110111101110, 25'b0000000000001001000001100, 25'b1111111111111101011010000, 25'b1111111111111100011110010, 25'b1111111111111100010010100, 25'b1111111111111111111001110, 25'b0000000000100010101100010, 25'b1111111111111111111111110, 25'b0000000000000000000000110, 25'b1111111111111110110011011, 25'b0000000000101000100111100, 25'b0000000000011000001010000, 25'b0000000000000100010110101, 25'b1111111111110011101010010, 25'b1111111111111110101111000, 25'b0000000000001000010110011, 25'b0000000000000111010111110},
{25'b0000000000000100010111001, 25'b0000000000000101000000000, 25'b1111111111111111111110101, 25'b0000000000000000000011011, 25'b1111111111000100000000101, 25'b0000000000000101100101101, 25'b0000000000000011001011101, 25'b1111111111111111111101111, 25'b0000000000000000000101110, 25'b1111111111101010010011110, 25'b1111111111111111111111111, 25'b0000000000000000000000010, 25'b1111111111101011011010101, 25'b0000000000000000000010000, 25'b0000000000000000000010101, 25'b0000000000000000000010111, 25'b0000000000000000000000011, 25'b1111111111010010011101100, 25'b0000000000000001001110001, 25'b1111111111111111111011110, 25'b1111111111111111111100110, 25'b0000000000000000000001011, 25'b0000000000010000100000100, 25'b1111111111111111111111010, 25'b0000000000000000000001001, 25'b0000000000111010010110101, 25'b0000000000101011100010101, 25'b0000000000000000000001100, 25'b0000000000000000000001011, 25'b1111111111100010000110110, 25'b0000000000000000000011001, 25'b1111111111111111111111011},
{25'b0000000000001001101100110, 25'b0000000000000110110000001, 25'b0000000000100000011001100, 25'b1111111111100000001110001, 25'b0000000000010000111100001, 25'b0000000000001111001100101, 25'b0000000000000000110011010, 25'b0000000000011000100011100, 25'b0000000000000001100001100, 25'b1111111111111110011101111, 25'b0000000000000100110001110, 25'b0000000000000000101111100, 25'b1111111111111111111011101, 25'b0000000000001111011100001, 25'b1111111111111111010010000, 25'b1111111111111010111011111, 25'b0000000000000000000101111, 25'b0000000000000100000100101, 25'b1111111111111001110101001, 25'b0000000000001100101000111, 25'b0000000000000100001010010, 25'b1111111110110101101101000, 25'b1111111111110001010110101, 25'b0000000000001011101100100, 25'b1111111111111111111111111, 25'b1111111110111111010111100, 25'b1111111111101111110110111, 25'b1111111111111101000011011, 25'b1111111111111111111010100, 25'b1111111111111000101100001, 25'b0000000000000000000000011, 25'b1111111111111010111100000},
{25'b0000000000000000001111000, 25'b1111111111111111111111001, 25'b1111111111110100010010101, 25'b1111111111101010011101100, 25'b0000000000000101010111111, 25'b0000000000000000000001110, 25'b0000000000001100001100111, 25'b1111111111111111010001001, 25'b0000000000011111111100101, 25'b1111111111111111011111000, 25'b0000000000000000000001000, 25'b1111111111010100000010100, 25'b1111111111111111111100111, 25'b0000000000010000000111110, 25'b1111111111111111111110011, 25'b1111111111011110101001000, 25'b0000000000000000000000100, 25'b1111111111111110100011010, 25'b0000000000100001101001111, 25'b1111111111111111111111101, 25'b1111111111001000000111110, 25'b1111111111111111111111000, 25'b0000000000100001000001110, 25'b1111111111111111111111011, 25'b1111111111111111111111010, 25'b0000000000010001110001111, 25'b1111111111110011111111011, 25'b0000000000001000110110101, 25'b0000000000000000000010000, 25'b1111111111100110001101110, 25'b0000000000000000000000111, 25'b0000000000000000010100001},
{25'b1111111111100100010101000, 25'b0000000000000000001001100, 25'b0000000000000000000100011, 25'b1111111111111111001110111, 25'b0000000000111111011101010, 25'b1111111111110000000110110, 25'b1111111111111111010010011, 25'b1111111111111111000100000, 25'b1111111111111010010001101, 25'b1111111111111001100011010, 25'b0000000000001000010110000, 25'b0000000000010001000000011, 25'b1111111111111011010010101, 25'b0000000000011111111100001, 25'b0000000000000000000001011, 25'b1111111111111111111101000, 25'b1111111111011011101000111, 25'b1111111111111111111011011, 25'b0000000000000000000011110, 25'b1111111111110101110011111, 25'b0000000000000000010001001, 25'b0000000000000100110001110, 25'b0000000000000001101101101, 25'b1111111111111110110101001, 25'b1111111111111001100000000, 25'b1111111111100110000010001, 25'b1111111111011010001000101, 25'b0000000000000000000010000, 25'b1111111111110001100000010, 25'b0000000000000101000110000, 25'b1111111111111111111101100, 25'b0000000000001001101011100},
{25'b1111111111001011000111011, 25'b1111111111101011111110110, 25'b1111111111101100000000101, 25'b0000000000000000000000110, 25'b0000000001001001000111110, 25'b1111111111100011100001000, 25'b0000000000000000000000100, 25'b1111111111111001000100010, 25'b1111111111001011100010110, 25'b0000000000010001101110111, 25'b1111111111111111111111111, 25'b0000000001001000100110001, 25'b0000000000000000000011101, 25'b1111111111111001111011100, 25'b1111111111111111111110000, 25'b0000000000000100000011101, 25'b1111111111111101100111110, 25'b0000000000000000000011100, 25'b1111111111111010000011000, 25'b0000000000111111011010011, 25'b0000000000000100111101101, 25'b1111111111111010101010011, 25'b0000000000001110000001010, 25'b1111111111111111111101101, 25'b1111111111111111111111101, 25'b1111111111110011100011111, 25'b1111111111111010000000011, 25'b1111111111000100000111010, 25'b1111111111101101100001000, 25'b1111111111111111111111101, 25'b1111111111111111110111100, 25'b1111111111111000011111101},
{25'b0000000000011100111010100, 25'b1111111110011001101010011, 25'b1111111110100011010001110, 25'b1111111111101010001110010, 25'b0000000001010101101011011, 25'b1111111111111111111111101, 25'b1111111111010011101000010, 25'b0000000000100001111001110, 25'b0000000000000111100110001, 25'b0000000000000000000111010, 25'b0000000000011010101011101, 25'b1111111111011101010000100, 25'b0000000000000000000111001, 25'b0000000000000000100011001, 25'b1111111111111011111111111, 25'b0000000000000010010011110, 25'b1111111111110010101101111, 25'b1111111110001010000011011, 25'b0000000000010101011110111, 25'b0000000000101100001001000, 25'b0000000000100001111100000, 25'b0000000000000000010101101, 25'b0000000000000011101110000, 25'b1111111111001100011011101, 25'b1111111110101111000000110, 25'b1111111111111111010111101, 25'b1111111111011001101000000, 25'b1111111111000101011001011, 25'b1111111111100111000011011, 25'b1111111110001111101111100, 25'b0000000000110101101010000, 25'b0000000000110110111100100},
{25'b0000000000000000000010000, 25'b0000000000000000000101001, 25'b0000000000000000010010011, 25'b0000000000000000000001101, 25'b0000000000100001001001010, 25'b1111111111101000000100010, 25'b0000000000000010010010000, 25'b0000000000001001010101110, 25'b1111111111010011010101001, 25'b0000000000000100101100111, 25'b1111111111111111011011001, 25'b1111111111111111111000010, 25'b1111111111111111111110100, 25'b0000000000011110101010111, 25'b0000000000000110101001001, 25'b0000000000000010110010000, 25'b0000000000000111111010011, 25'b0000000000101010101010001, 25'b1111111111100100000010100, 25'b0000000000000000000001000, 25'b1111111111101010111110011, 25'b1111111111111111111101101, 25'b0000000000101000010001111, 25'b0000000000000001000010110, 25'b1111111111111111101001000, 25'b1111111110111000001011100, 25'b1111111111111110110101000, 25'b1111111111101100001111101, 25'b1111111111111000001100110, 25'b0000000000000000011101001, 25'b0000000000010001010010100, 25'b0000000000001101010001100},
{25'b1111111111111010011101101, 25'b0000000000010001001001001, 25'b1111111111011001000111001, 25'b0000000000000010101001100, 25'b0000000000011000110010011, 25'b1111111111111010111100000, 25'b1111111111111111011010001, 25'b0000000000010100111001111, 25'b0000000000000000000010010, 25'b1111111111111111111110011, 25'b1111111111110111101000010, 25'b0000000000000000000000010, 25'b0000000000000000000011001, 25'b1111111111111011100111110, 25'b1111111111110000011011001, 25'b1111111111110111100000110, 25'b1111111111111000110010010, 25'b1111111111110111111101010, 25'b1111111111110001111100101, 25'b0000000000000000000001000, 25'b1111111111111111111101101, 25'b1111111111111010010001111, 25'b1111111111110111011110001, 25'b0000000000110010111010110, 25'b0000000000000000000000010, 25'b1111111111010001111011001, 25'b1111111111111110111010110, 25'b0000000000001111110001011, 25'b0000000000000000000011100, 25'b0000000000000000000000000, 25'b0000000000100000001000000, 25'b1111111111111111111100101},
{25'b1111111111111111111111001, 25'b0000000000000000100001101, 25'b1111111111111111111101001, 25'b1111111111101100000000001, 25'b1111111110010001111000011, 25'b0000000000000000000111100, 25'b0000000000000000000010101, 25'b1111111111111111001010110, 25'b1111111110110011010000101, 25'b0000000000001010011100011, 25'b1111111111110011011100110, 25'b1111111111111111111111100, 25'b0000000000000000000011111, 25'b1111111111010000101001100, 25'b1111111111111010001001000, 25'b1111111111111111111101110, 25'b0000000000000000001011001, 25'b0000000000000001000011110, 25'b0000000000000100101001011, 25'b0000000000101100001100011, 25'b1111111111110000101100000, 25'b1111111111011001101110100, 25'b0000000000000000000000111, 25'b1111111111011110111111101, 25'b1111111111110011010111110, 25'b1111111111100010011000111, 25'b1111111111111111000011100, 25'b1111111111111110011001100, 25'b1111111111111101101011010, 25'b1111111111000011101100101, 25'b1111111111111011101000111, 25'b0000000000011111000000101},
{25'b0000000000001110011111101, 25'b0000000000011100000011101, 25'b1111111111111111101111110, 25'b0000000000010100011001001, 25'b1111111111100101000000001, 25'b1111111111110000000100100, 25'b0000000000001100001111011, 25'b0000000000001000110010101, 25'b1111111111111001111110100, 25'b1111111111111111111111000, 25'b1111111111111111111111000, 25'b1111111111111111111110010, 25'b1111111111111111111101100, 25'b1111111111010110111111110, 25'b1111111111111111111111011, 25'b0000000000010010011101100, 25'b1111111111110001010111100, 25'b0000000000000100011101011, 25'b1111111111111111110101001, 25'b1111111111111111110111101, 25'b0000000000011010100011000, 25'b1111111111010110001000100, 25'b0000000000100011111100101, 25'b0000000000000110000101010, 25'b0000000000000000000010001, 25'b0000000000011011000111111, 25'b0000000000000000011010000, 25'b1111111111111011011000010, 25'b1111111111001111010011000, 25'b1111111111110001111111110, 25'b1111111111101010001101011, 25'b0000000000010110101110101},
{25'b0000000000000000000000010, 25'b0000000000000000111011000, 25'b1111111111010001001010111, 25'b1111111111111111101100010, 25'b0000000000011010011101100, 25'b1111111111101101111000010, 25'b1111111111111110011101010, 25'b1111111111111111111111011, 25'b0000000000000010100110111, 25'b0000000000000000000000011, 25'b0000000000000000000000010, 25'b1111111111100101111010100, 25'b0000000000001100010010100, 25'b0000000000000000110001101, 25'b0000000000000000000001010, 25'b0000000000000100110010110, 25'b1111111111111111111101011, 25'b1111111111101100111101110, 25'b0000000000000010010010101, 25'b0000000000000000000001011, 25'b1111111111111011100110111, 25'b1111111111111101001100100, 25'b0000000000100101111011011, 25'b1111111111111111111111010, 25'b0000000000000000000000100, 25'b1111111111011010100010100, 25'b1111111111010110001010100, 25'b0000000000011110111001111, 25'b1111111111111111110101110, 25'b1111111111111111111101001, 25'b0000000000000011100010111, 25'b0000000000100100001011100},
{25'b1111111111010100011000100, 25'b1111111111111111111111100, 25'b1111111111100100110001101, 25'b0000000000000000100011000, 25'b1111111111010010110001011, 25'b0000000000000000000000000, 25'b1111111111111111111101111, 25'b1111111111110111101000100, 25'b1111111110111011110111100, 25'b1111111111111100101101010, 25'b0000000000000000000000110, 25'b1111111111111110111100001, 25'b1111111111111111111101010, 25'b0000000000000000000000110, 25'b1111111111111110111001111, 25'b1111111111111001101000101, 25'b1111111111101101000111110, 25'b1111111111110011110010110, 25'b0000000000001000011110100, 25'b1111111111111111101100100, 25'b1111111111111100110000111, 25'b0000000000000000000000101, 25'b0000000000101011000110000, 25'b1111111111111111111110111, 25'b0000000000010011001000010, 25'b0000000000001011101111010, 25'b1111111111101110011000110, 25'b0000000000011011010011010, 25'b1111111111111010001001010, 25'b0000000000000000000000011, 25'b1111111111111111110110110, 25'b0000000001001010100000001},
{25'b1111111111010111110011111, 25'b0000000000000011110011100, 25'b0000000000000110011111000, 25'b1111111111111100011010000, 25'b0000000000011111010000110, 25'b1111111111011001010100000, 25'b1111111111111111000110110, 25'b0000000000100001111111111, 25'b0000000000010100011001000, 25'b0000000000000001001011100, 25'b1111111111111111111111001, 25'b1111111111110111001111100, 25'b1111111111110100100011001, 25'b1111111111110111101110001, 25'b1111111111111001101001011, 25'b0000000000001011100011001, 25'b1111111111111111111111000, 25'b0000000000000001000010011, 25'b0000000000010010000101111, 25'b0000000000000000000000110, 25'b0000000000000000000001000, 25'b0000000000000001111010100, 25'b0000000000100000010000100, 25'b0000000000000101110110100, 25'b0000000000000000110110110, 25'b1111111111110010001110101, 25'b1111111111111111111111010, 25'b0000000000000000000000010, 25'b1111111111111110001100000, 25'b1111111111111110011101001, 25'b1111111111111111111101100, 25'b0000000000001000101001101},
{25'b1111111111111111111110101, 25'b0000000000000000011111101, 25'b1111111111100100110111011, 25'b1111111111110110011101101, 25'b0000000000100100000111100, 25'b1111111111111111111101010, 25'b1111111111110110000110000, 25'b0000000000011111010010111, 25'b1111111111111001001110010, 25'b0000000000100101010101010, 25'b0000000000001010111100110, 25'b1111111111110000100111100, 25'b0000000000000000000100101, 25'b0000000000000000011100111, 25'b1111111111111110000111111, 25'b0000000000000010101110001, 25'b1111111111110110001000110, 25'b1111111111011110010011001, 25'b0000000000100011100101000, 25'b0000000000010011111000100, 25'b0000000001010001001111100, 25'b0000000000011001101100001, 25'b0000000000011111110000011, 25'b1111111111111111111110001, 25'b0000000000000000000000010, 25'b0000000000000000000000011, 25'b0000000000000111010101111, 25'b0000000000001010001001010, 25'b1111111111001010010000000, 25'b1111111111111111111110011, 25'b1111111111111111010110001, 25'b1111111111111111001010010},
{25'b0000000000000000000100010, 25'b1111111111110100110010010, 25'b1111111111110010101111111, 25'b0000000000000000000000100, 25'b1111111111100000110100000, 25'b0000000000000000000000101, 25'b0000000000011000100000011, 25'b0000000000001101111110010, 25'b0000000000000110110011001, 25'b1111111111110011010111010, 25'b0000000000000000000000101, 25'b1111111111111111111111101, 25'b1111111111111111111110001, 25'b1111111111111111111110101, 25'b1111111111111010100010101, 25'b0000000000011001110111001, 25'b1111111111111111111111101, 25'b1111111111111111111011111, 25'b1111111111011001010011011, 25'b0000000000000000000001100, 25'b1111111111100111010111111, 25'b1111111111111111110111111, 25'b0000000000000000000001100, 25'b1111111111111111011110011, 25'b0000000000000001111011100, 25'b0000000000000010001111000, 25'b0000000000000011100100111, 25'b0000000000010001101101110, 25'b1111111111110111101011100, 25'b1111111111111111000001011, 25'b1111111111000110100100110, 25'b0000000000001010000101110},
{25'b0000000000111000100011011, 25'b1111111111111110111000111, 25'b0000000000001000011110100, 25'b1111111111110010100110011, 25'b1111111111110101000100101, 25'b0000000000000100010001011, 25'b0000000000010100100000101, 25'b0000000000000000000000110, 25'b0000000001000011011101011, 25'b0000000000000000000010101, 25'b1111111111111101010000101, 25'b0000000000000010011010110, 25'b0000000000001100000010101, 25'b1111111111111111101010110, 25'b0000000000000110110100001, 25'b0000000000001101001110100, 25'b1111111111111111011101000, 25'b1111111111000111000001011, 25'b1111111111111000110010000, 25'b1111111111111111110010100, 25'b0000000000001110111000101, 25'b0000000000000000001110000, 25'b1111111111111111111100001, 25'b0000000000001110011001100, 25'b0000000000000010010011001, 25'b1111111111011110010000101, 25'b1111111111110010110110110, 25'b0000000000010000111011010, 25'b1111111111111100011000101, 25'b0000000000100001000010011, 25'b1111111111111111110111001, 25'b1111111111101001000111111},
{25'b0000000000000001101010010, 25'b0000000000001101000010111, 25'b1111111111111111111111101, 25'b1111111111111011000010111, 25'b1111111111010010110100100, 25'b1111111111111111111100110, 25'b0000000000000101111001000, 25'b1111111111111010000111000, 25'b0000000000010101000111000, 25'b1111111111111011101000001, 25'b1111111111111111111001010, 25'b1111111111111011101110011, 25'b1111111111111111111110000, 25'b1111111111111011010000111, 25'b0000000000000000000000110, 25'b0000000000101000000100110, 25'b0000000000000000000000100, 25'b1111111111111111110010000, 25'b1111111111111111111110001, 25'b1111111111111111111110101, 25'b1111111111111111111110001, 25'b1111111111111111111100101, 25'b0000000000000100010111100, 25'b0000000000010000000111100, 25'b0000000000000000000000001, 25'b0000000000000000100010001, 25'b0000000000000100001001011, 25'b1111111111111111111011101, 25'b0000000000000000000000110, 25'b0000000000000010100111001, 25'b0000000000000000001100011, 25'b0000000000001100011001000},
{25'b1111111111011000011110000, 25'b0000000000010000101011010, 25'b0000000000000010010011010, 25'b1111111111110010100011111, 25'b1111111111001100111001001, 25'b1111111111111101101010000, 25'b0000000000001000100100110, 25'b1111111111001101001000010, 25'b0000000001000001011110110, 25'b0000000000001001001011000, 25'b0000000000000010000000001, 25'b0000000000001100000100010, 25'b0000000000000101101011011, 25'b0000000000000000000101101, 25'b0000000000110100001100111, 25'b1111111111110101001110111, 25'b0000000000000000101010101, 25'b0000000000000000000000111, 25'b1111111111111111001001001, 25'b0000000000000000011110111, 25'b1111111111001000101111000, 25'b0000000000000010001010111, 25'b0000000000010011100100101, 25'b0000000000000100110011111, 25'b0000000000000100100111110, 25'b1111111110101011111111101, 25'b1111111111010100010111110, 25'b1111111111100001001100100, 25'b0000000000000000010101111, 25'b1111111111111111110001100, 25'b0000000000101001101110000, 25'b1111111111100101110010110},
{25'b1111111111111110010110110, 25'b1111111111100111001000000, 25'b1111111111110010110001001, 25'b1111111111001011101100011, 25'b1111111111011110101100101, 25'b0000000000101011000010010, 25'b0000000000100111101010101, 25'b1111111111101010001110101, 25'b0000000000000101010100110, 25'b1111111111111011000010100, 25'b1111111111110011111110101, 25'b1111111111011111110100111, 25'b0000000000001101001100111, 25'b1111111111011011101000001, 25'b0000000000011000001010001, 25'b1111111111111111111101010, 25'b0000000000101010111111100, 25'b1111111111111111111111111, 25'b1111111111111111000000000, 25'b1111111111101110101011001, 25'b1111111111111010101011011, 25'b1111111111110111101111111, 25'b1111111111011110000000000, 25'b0000000000001010100010111, 25'b1111111111111111111111001, 25'b1111111111111111001100010, 25'b1111111111100010110010111, 25'b0000000000101000010011100, 25'b0000000000100011101110010, 25'b1111111111110100011011000, 25'b1111111110101111010010111, 25'b0000000000010010010010010},
{25'b0000000000000000000011001, 25'b1111111111111100101110101, 25'b1111111111111111111110010, 25'b1111111111110011100011110, 25'b0000000000000011101001011, 25'b0000000000000001001010110, 25'b0000000000001000111010111, 25'b0000000000000000101111010, 25'b0000000000001111000101110, 25'b1111111111111111111000011, 25'b0000000000000000000000000, 25'b0000000000001100001101110, 25'b0000000000000000001111001, 25'b0000000000000001100100001, 25'b1111111111101111000100000, 25'b1111111111110010001101110, 25'b0000000000000000000000101, 25'b0000000000010111010001000, 25'b0000000000000111010001100, 25'b0000000000010000000110001, 25'b1111111111111101111000101, 25'b1111111111101011100010101, 25'b1111111111111111111110100, 25'b0000000000001001100000101, 25'b1111111111111111111110111, 25'b0000000000000100001001010, 25'b1111111111111111011000100, 25'b0000000000001000101001010, 25'b0000000000000000000001110, 25'b0000000000001010101001011, 25'b1111111111001111011011011, 25'b1111111111111111111111011},
{25'b0000000000100111101111000, 25'b1111111111111110110110010, 25'b0000000000010011001100010, 25'b1111111111011000111011100, 25'b1111111111100111010010010, 25'b1111111111111111111111010, 25'b1111111111111111111110111, 25'b0000000000000011100000001, 25'b0000000000000000010011000, 25'b1111111111101111111000011, 25'b0000000000000000000000001, 25'b0000000000000000010000001, 25'b0000000000000000000000010, 25'b0000000000000000000010110, 25'b1111111111101111011110011, 25'b0000000000010010010000011, 25'b1111111111111111110010111, 25'b1111111111111100000011000, 25'b0000000000000000000001010, 25'b0000000000001111010111011, 25'b1111111111100110010011001, 25'b0000000000001110110111111, 25'b0000000000010001111011110, 25'b0000000000010000100000100, 25'b1111111111111111111111101, 25'b0000000001000110100101110, 25'b1111111111101100011001110, 25'b0000000000101110100001001, 25'b1111111111111001011010000, 25'b1111111111010001110101101, 25'b1111111111101001110011110, 25'b0000000000010001110110001},
{25'b1111111110111010011110111, 25'b1111111111111100100101010, 25'b1111111111101100010010011, 25'b1111111111111111111111101, 25'b0000000000100001011000011, 25'b1111111111101001001001101, 25'b1111111111111000010101010, 25'b0000000000011110011111110, 25'b0000000000001100000110111, 25'b1111111111100001100010100, 25'b0000000000000000000001010, 25'b1111111111111100011001100, 25'b1111111111111110101111110, 25'b0000000000010001100110110, 25'b1111111111100000100011100, 25'b1111111111111110100100011, 25'b0000000000000000000000100, 25'b1111111111111111111010110, 25'b1111111111111101111100101, 25'b0000000000000000000001000, 25'b1111111111100111101010110, 25'b1111111111111111111110011, 25'b0000000000000000000000101, 25'b1111111111010101111110011, 25'b0000000000001000111111001, 25'b0000000001001111010101111, 25'b0000000000101100010001001, 25'b1111111111111011011010101, 25'b1111111111101011011100101, 25'b1111111111000110100100110, 25'b0000000000000000000010110, 25'b1111111111111001110000010},
{25'b0000000000000010101111100, 25'b0000000000011011010110111, 25'b0000000000000010101110010, 25'b1111111111101100101010001, 25'b0000000000000000100101110, 25'b1111111111111100101111110, 25'b0000000000000000000001101, 25'b0000000000011010101011110, 25'b0000000000011011100000110, 25'b1111111111101110111001010, 25'b0000000000010001111111000, 25'b0000000000000011000100111, 25'b1111111111111111111111011, 25'b1111111111111110001011011, 25'b1111111111101011101011010, 25'b0000000000100000011000001, 25'b1111111111111010100100110, 25'b1111111111010110101001001, 25'b0000000000001110101000110, 25'b1111111111111111111110110, 25'b1111111111111111111110010, 25'b0000000000001110111101011, 25'b1111111111110110011111001, 25'b1111111111111111011000100, 25'b1111111111111001011001011, 25'b0000000000001011010010001, 25'b1111111111101110000010110, 25'b0000000000010001001010111, 25'b1111111111010001011100001, 25'b0000000000001010010011010, 25'b1111111111111111111100011, 25'b0000000000010100000011011},
{25'b1111111111111010100000101, 25'b0000000000000000000100111, 25'b0000000000001011011001011, 25'b0000000000000000000000111, 25'b1111111111111000001100001, 25'b1111111111111111101000101, 25'b0000000000001101001000111, 25'b1111111111111111111111101, 25'b0000000000000000000010000, 25'b0000000000000000101001101, 25'b0000000000000000000001011, 25'b0000000000000010100011010, 25'b1111111111110010011001011, 25'b0000000000000001010101011, 25'b0000000000001110001011011, 25'b0000000000000101111110110, 25'b0000000000001101100000110, 25'b1111111111111111111011110, 25'b1111111111111111110101001, 25'b0000000000010000011000100, 25'b0000000000011111101010110, 25'b1111111111110011011110110, 25'b0000000000000000000000100, 25'b1111111111111111101111010, 25'b0000000000000001011101101, 25'b1111111111000100111111101, 25'b1111111111111111111001011, 25'b1111111111110110111100010, 25'b1111111111111111111110010, 25'b0000000001001000010001000, 25'b0000000000000000000010010, 25'b1111111111100101101001010},
{25'b1111111111111100100100001, 25'b1111111111110000101110011, 25'b1111111111111110110111111, 25'b0000000000000000111001100, 25'b0000000000001011100111010, 25'b1111111111111111111111001, 25'b0000000000000000000010000, 25'b1111111111111101000010100, 25'b0000000000001001000011000, 25'b1111111111111110111100111, 25'b0000000000000000000001010, 25'b0000000000000100000011100, 25'b0000000000100101110000111, 25'b1111111111110010111100101, 25'b0000000000000001100111010, 25'b1111111110010011011011011, 25'b1111111111111110100100110, 25'b1111111111111000010000100, 25'b0000000000000001000001100, 25'b1111111111111001100111001, 25'b0000000000001011110001110, 25'b1111111111100011010100000, 25'b0000000000001110100111010, 25'b0000000000001101011111101, 25'b1111111111111110010100101, 25'b1111111110100100111111010, 25'b1111111111100010101111111, 25'b1111111111111101001101001, 25'b1111111111111101101001110, 25'b0000000000110001111111011, 25'b1111111111111111010000100, 25'b0000000000010011101110100},
{25'b0000000000000110000000111, 25'b0000000000000000000001011, 25'b0000000000010110010010111, 25'b1111111111110001011111000, 25'b1111111111110111001100111, 25'b0000000000011110011100110, 25'b1111111111101011100010010, 25'b0000000000000111010111000, 25'b1111111111011000011001011, 25'b0000000000000001000111111, 25'b0000000000000010001001011, 25'b1111111111110101010001000, 25'b0000000000000000000100011, 25'b0000000000000000000000000, 25'b1111111111100111111101000, 25'b0000000000110111010111000, 25'b1111111111100000011010110, 25'b1111111111111110011110100, 25'b0000000000001111001101101, 25'b1111111111111111111110111, 25'b0000000000001000110111110, 25'b1111111111000010101011001, 25'b0000000000101000000101100, 25'b1111111111111111111111100, 25'b1111111111110000001001101, 25'b0000000000111110000010011, 25'b0000000000010010101100100, 25'b1111111111101011110011100, 25'b1111111111101110110011000, 25'b1111111110111011001111110, 25'b1111111111111110101100101, 25'b0000000000000010000010001},
{25'b1111111111111111111111110, 25'b0000000000000000110101111, 25'b1111111111111011100011011, 25'b1111111111011101101100111, 25'b1111111111111111111101011, 25'b1111111111001101110001011, 25'b0000000000000000000010011, 25'b0000000000100110110111001, 25'b0000000000011111010001010, 25'b0000000000000010011010110, 25'b0000000000000000000000001, 25'b1111111111110001111001110, 25'b0000000000101010100000110, 25'b1111111111111111111111110, 25'b1111111111111111111101100, 25'b1111111111111111111100101, 25'b0000000000110111100010110, 25'b0000000000000000001101000, 25'b1111111111111010111010100, 25'b1111111111111001011101111, 25'b1111111111010110110011011, 25'b0000000000010000110110000, 25'b0000000000000000000000001, 25'b0000000000000000000000011, 25'b0000000000000100000011001, 25'b1111111111110110111001011, 25'b1111111111000101000010111, 25'b0000000000100011010100010, 25'b1111111111000111001111110, 25'b0000000000000110100010111, 25'b1111111111110101111001100, 25'b0000000000000000000000001},
{25'b0000000000000111110110001, 25'b0000000000010111110111011, 25'b0000000000000001001111000, 25'b1111111111111111100111101, 25'b1111111111000101001110000, 25'b0000000000000000000111100, 25'b1111111111111111111111101, 25'b0000000000011111000000111, 25'b0000000000100011011101100, 25'b1111111111111111111110101, 25'b1111111111111111111110111, 25'b1111111111111111110110000, 25'b0000000000000000000001011, 25'b0000000000000000010000111, 25'b0000000000000000000000000, 25'b0000000000000000000001110, 25'b0000000000000000000011101, 25'b1111111111111111111010111, 25'b0000000000010101110000001, 25'b1111111111110010110100101, 25'b1111111111001000101101010, 25'b1111111111111011110000100, 25'b1111111111110011010110000, 25'b1111111111110011111111100, 25'b1111111111110111001000111, 25'b1111111111111111111000100, 25'b1111111111110111111100110, 25'b1111111111111101001100101, 25'b1111111111111110101010111, 25'b0000000000010010000110110, 25'b1111111111111111111101011, 25'b0000000000111011010100101}
};
localparam logic signed [24:0] bias [32] = '{
25'b0000000010111100101101010,
25'b0000000001011000100000101,
25'b0000000010111000011001110,
25'b0000000010110100001110110,
25'b0000000001111110010001010,
25'b0000000001101110100010110,
25'b1111111110110001001111000,
25'b0000000000111101111100010,
25'b0000000000111110001111101,
25'b0000000000101111100100011,
25'b0000000000111010110111100,
25'b0000000010100110011000001,
25'b1111111101111101111000101,
25'b1111111111010010111000011,
25'b0000000000111001000100001,
25'b1111111111110001101010100,
25'b1111111111110111011001110,
25'b0000000000000000101000000,
25'b0000000000011000111010111,
25'b1111111110011100001100111,
25'b0000000001011101010001111,
25'b0000000011011011100000010,
25'b1111111100110011100100100,
25'b0000000000001001011101101,
25'b0000000000101001010010011,
25'b0000000001101100001101000,
25'b0000000001110011000001010,
25'b0000000000100000101000000,
25'b0000000001111100100111100,
25'b0000000010010000001001110,
25'b0000000000111001010011011,
25'b1111111011010000111100101
};
endpackage