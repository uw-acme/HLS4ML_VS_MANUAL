// Width: 11
// NFRAC: 5
package dense_1_11_5;

localparam logic signed [10:0] weights [16][64] = '{ 
{11'b00000001000, 11'b11111101011, 11'b11111111010, 11'b11111111000, 11'b11111110011, 11'b00000000011, 11'b11111011110, 11'b00000000000, 11'b00000000001, 11'b00000001000, 11'b00000000000, 11'b11111110011, 11'b11111111111, 11'b00000000110, 11'b00000000001, 11'b11111110111, 11'b00000000111, 11'b00000000001, 11'b00000000000, 11'b11111111111, 11'b00000001100, 11'b11111110101, 11'b11111111111, 11'b00000001111, 11'b11111110101, 11'b11111101010, 11'b11111110111, 11'b11111111001, 11'b11111111100, 11'b11111111111, 11'b00000000001, 11'b00000000111, 11'b00000000110, 11'b11111111111, 11'b00000000000, 11'b00000001001, 11'b11111111111, 11'b11111110111, 11'b00000000000, 11'b00000000110, 11'b11111111111, 11'b00000001000, 11'b11111110111, 11'b00000011101, 11'b11111111111, 11'b00000001110, 11'b00000000000, 11'b00000000101, 11'b00000000110, 11'b11111111111, 11'b00000000000, 11'b00000000101, 11'b00000000110, 11'b00000000010, 11'b11111111100, 11'b11111110110, 11'b00000010001, 11'b11111110000, 11'b00000001110, 11'b11111110100, 11'b00000011001, 11'b11111111111, 11'b00000000000, 11'b00000000010}, 
{11'b00000000000, 11'b11111110101, 11'b11111111011, 11'b11111110111, 11'b11111110101, 11'b00000000011, 11'b11111100111, 11'b11111111111, 11'b11111111000, 11'b00000000101, 11'b00000000000, 11'b11111111101, 11'b00000000110, 11'b00000000000, 11'b11111111111, 11'b00000000110, 11'b11111111111, 11'b00000000000, 11'b11111111010, 11'b11111110111, 11'b00000001110, 11'b11111111101, 11'b00000000001, 11'b00000010110, 11'b00000001000, 11'b11111111000, 11'b11111111000, 11'b11111111111, 11'b11111111100, 11'b11111110011, 11'b11111111110, 11'b00000001110, 11'b00000001000, 11'b00000010001, 11'b00000010100, 11'b00000000001, 11'b11111111100, 11'b11111110010, 11'b00000000001, 11'b00000000110, 11'b00000000000, 11'b00000000110, 11'b11111111001, 11'b00000001000, 11'b00000000101, 11'b00000000001, 11'b11111110101, 11'b00000000010, 11'b00000001000, 11'b00000000000, 11'b00000000000, 11'b00000100101, 11'b11111111101, 11'b11111111100, 11'b11111111110, 11'b11111111111, 11'b00000001000, 11'b11111110100, 11'b00000011111, 11'b00000000000, 11'b00000010000, 11'b00000000111, 11'b00000011010, 11'b00000000100}, 
{11'b11111111111, 11'b00000000000, 11'b11111111101, 11'b11111111010, 11'b11111111010, 11'b00000000001, 11'b00000101111, 11'b11111111111, 11'b11111010111, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b11111111000, 11'b00000000000, 11'b11111111111, 11'b00000000101, 11'b00000011100, 11'b11111111111, 11'b00000000010, 11'b00000000000, 11'b00000001101, 11'b11111101000, 11'b00000010010, 11'b11111101001, 11'b00000011110, 11'b11111110100, 11'b11111111000, 11'b11111101001, 11'b00000101000, 11'b00000001000, 11'b00000000000, 11'b00000010000, 11'b00000100000, 11'b11111011001, 11'b11111111100, 11'b00000000001, 11'b11111111000, 11'b00000011100, 11'b11111111110, 11'b00000001010, 11'b00000001010, 11'b00000001011, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b00000000101, 11'b11111110111, 11'b11111111010, 11'b11111111111, 11'b00000001100, 11'b11111111010, 11'b00000000100, 11'b11111111111, 11'b00000000100, 11'b11111111010, 11'b11111111111, 11'b11111110110, 11'b11111101010, 11'b11111111111, 11'b00000000000, 11'b00000110001, 11'b00000000000, 11'b11111111111, 11'b11111110110}, 
{11'b11111110001, 11'b11111110100, 11'b11111101001, 11'b00000001001, 11'b11111110101, 11'b11111010100, 11'b11111111100, 11'b11111110110, 11'b00000000111, 11'b11111111111, 11'b00000101000, 11'b11111111100, 11'b11111100110, 11'b00000010010, 11'b00000000000, 11'b11111111111, 11'b11111110001, 11'b11111111111, 11'b00000000000, 11'b11111111000, 11'b11111011011, 11'b11111111100, 11'b11111101001, 11'b00000000110, 11'b11111110011, 11'b11111100010, 11'b00000001010, 11'b00000010111, 11'b00000101001, 11'b11111110001, 11'b11111101101, 11'b00000000010, 11'b00000010000, 11'b11111100101, 11'b11111110101, 11'b00000000000, 11'b11111101000, 11'b00000000111, 11'b11111110001, 11'b00000000011, 11'b00000001110, 11'b00000000101, 11'b00000000000, 11'b00000000000, 11'b00000010001, 11'b11111111001, 11'b11111111111, 11'b11111110100, 11'b11111111111, 11'b11111111100, 11'b11111101100, 11'b00000000010, 11'b11111111111, 11'b00000000110, 11'b00000001010, 11'b00000010100, 11'b11111100001, 11'b11111100010, 11'b11111101001, 11'b00000011011, 11'b00000110111, 11'b11111100011, 11'b11111111110, 11'b00000001101}, 
{11'b00000001010, 11'b11111101100, 11'b11111110111, 11'b11111111111, 11'b11111111011, 11'b00000001010, 11'b00000000110, 11'b11111111111, 11'b11111101100, 11'b11111111000, 11'b11111110100, 11'b00000000001, 11'b00000000000, 11'b00000000000, 11'b11111111110, 11'b00000001011, 11'b00000000100, 11'b11111110011, 11'b00000000000, 11'b00000000000, 11'b00000000110, 11'b11111111100, 11'b00000000010, 11'b11111111111, 11'b00000100010, 11'b11111111010, 11'b11111110111, 11'b11111110011, 11'b00000000000, 11'b00000000101, 11'b00000000011, 11'b00000001000, 11'b11111111111, 11'b00000000010, 11'b00000000100, 11'b11111111111, 11'b00000000000, 11'b00000011100, 11'b11111110110, 11'b11111111101, 11'b00000001101, 11'b00000000111, 11'b11111110000, 11'b00000000000, 11'b11111011101, 11'b11111111111, 11'b11111111100, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b00000000110, 11'b11111111111, 11'b00000001010, 11'b11111111001, 11'b11111101000, 11'b11111110001, 11'b11111101111, 11'b11111101100, 11'b00000010111, 11'b00000101011, 11'b00000011001, 11'b00000000011, 11'b11111111111}, 
{11'b11111110001, 11'b11111101011, 11'b00000000000, 11'b00000001001, 11'b00000001001, 11'b11111111001, 11'b00000010010, 11'b11111111111, 11'b00000000111, 11'b11111111111, 11'b11111111111, 11'b11111111101, 11'b11111111010, 11'b00000010010, 11'b11111111101, 11'b00000000000, 11'b11111101100, 11'b11111110100, 11'b00000000000, 11'b11111111111, 11'b11111111110, 11'b11111110101, 11'b11111110101, 11'b00000001110, 11'b11111110101, 11'b11111111111, 11'b00000001000, 11'b11111111101, 11'b11111100010, 11'b11111111111, 11'b11111111101, 11'b11111111111, 11'b11111111111, 11'b00000000001, 11'b00000000100, 11'b00000001011, 11'b00000000000, 11'b11111111100, 11'b11111110111, 11'b11111111111, 11'b11111111010, 11'b11111101111, 11'b00000001100, 11'b00000000000, 11'b00000010011, 11'b00000000000, 11'b11111111111, 11'b00000000011, 11'b11111110010, 11'b00000000111, 11'b00000000000, 11'b11111111100, 11'b11111110100, 11'b00000001100, 11'b11111111111, 11'b00000001011, 11'b00000000110, 11'b00000000110, 11'b11111111111, 11'b11111111111, 11'b11111100110, 11'b11111111011, 11'b11111111110, 11'b11111111111}, 
{11'b11111110110, 11'b11111110101, 11'b11111110010, 11'b11111111101, 11'b11111111011, 11'b00000000011, 11'b11111101001, 11'b11111111011, 11'b11111111000, 11'b11111111111, 11'b11111110110, 11'b00000001011, 11'b00000000001, 11'b00000000100, 11'b00000001001, 11'b00000000000, 11'b00000011001, 11'b00000000010, 11'b00000000111, 11'b00000001000, 11'b11111111010, 11'b00000001011, 11'b11111111000, 11'b11111101111, 11'b00000000101, 11'b00000010000, 11'b11111111111, 11'b00000000001, 11'b11111100001, 11'b00000001001, 11'b00000001000, 11'b11111110100, 11'b00000001111, 11'b00000010101, 11'b00000000000, 11'b00000001010, 11'b11111111111, 11'b00000001001, 11'b00000000110, 11'b00000000000, 11'b11111111100, 11'b11111110100, 11'b00000000100, 11'b00000001111, 11'b00000010000, 11'b11111111010, 11'b11111111101, 11'b11111111001, 11'b11111111011, 11'b00000000011, 11'b00000000000, 11'b00000000001, 11'b00000000000, 11'b00000000101, 11'b11111111010, 11'b00000011000, 11'b00000001011, 11'b11111111111, 11'b00000001100, 11'b00000000110, 11'b11111001011, 11'b11111101101, 11'b11111111010, 11'b11111111111}, 
{11'b00000000000, 11'b00000000111, 11'b11111111111, 11'b11111111111, 11'b11111110101, 11'b11111111111, 11'b11111110111, 11'b00000000000, 11'b00000000000, 11'b00000001100, 11'b00000000000, 11'b11111110011, 11'b11111111101, 11'b00000000000, 11'b11111111110, 11'b11111110001, 11'b11111100100, 11'b11111111111, 11'b11111101100, 11'b11111110001, 11'b11111110011, 11'b00000001011, 11'b00000000001, 11'b11111111011, 11'b11111110010, 11'b00000000100, 11'b00000000000, 11'b00000001111, 11'b00000011001, 11'b11111111110, 11'b00000000000, 11'b00000000111, 11'b11111101010, 11'b11111110100, 11'b00000000001, 11'b00000000010, 11'b11111110111, 11'b00000000111, 11'b00000000100, 11'b11111111011, 11'b11111110010, 11'b11111111110, 11'b00000000001, 11'b11111111010, 11'b00000000001, 11'b00000000111, 11'b11111111100, 11'b00000000000, 11'b00000000000, 11'b11111111001, 11'b11111110011, 11'b00000001101, 11'b00000000100, 11'b11111111010, 11'b00000000100, 11'b11111111110, 11'b11111110000, 11'b11111111011, 11'b11111111110, 11'b11111111101, 11'b00000011010, 11'b00000000110, 11'b11111111110, 11'b11111111111}, 
{11'b00000000000, 11'b00000010010, 11'b11111101101, 11'b11111111000, 11'b00000001010, 11'b11111111001, 11'b00000100110, 11'b11111110110, 11'b11111111111, 11'b00000001001, 11'b00000001000, 11'b11111111111, 11'b11111111110, 11'b11111110000, 11'b00000001001, 11'b00000000101, 11'b11111111001, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b00000001000, 11'b11111110001, 11'b00000001100, 11'b00000010011, 11'b11111111101, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b00000010111, 11'b00000000000, 11'b11111110111, 11'b00000000000, 11'b00000001100, 11'b11111100110, 11'b11111101110, 11'b00000000110, 11'b00000000100, 11'b11111101101, 11'b11111111001, 11'b11111111001, 11'b00000001100, 11'b00000001100, 11'b00000000000, 11'b11111110111, 11'b00000000000, 11'b00000001100, 11'b11111111110, 11'b11111111111, 11'b00000000000, 11'b00000000111, 11'b11111111110, 11'b11111111001, 11'b00000001011, 11'b11111111001, 11'b00000001000, 11'b00000010010, 11'b00000000001, 11'b00000001000, 11'b11111110011, 11'b11111110100, 11'b00000011010, 11'b11111111011, 11'b00000000001, 11'b11111111101}, 
{11'b00000000000, 11'b11111110001, 11'b00000001011, 11'b11111110110, 11'b11111111111, 11'b00000000110, 11'b11111101101, 11'b00000000110, 11'b00000001111, 11'b00000000100, 11'b00000001011, 11'b00000001010, 11'b11111110110, 11'b11111111101, 11'b11111111110, 11'b00000000000, 11'b11111100001, 11'b00000001010, 11'b11111111110, 11'b00000000000, 11'b11111110100, 11'b00000000010, 11'b00000000100, 11'b11111111111, 11'b11111110001, 11'b11111111110, 11'b11111111101, 11'b00000100111, 11'b11111101010, 11'b00000000010, 11'b00000000011, 11'b11111111110, 11'b11111111000, 11'b00000000011, 11'b11111111101, 11'b11111111011, 11'b11111111010, 11'b11111111001, 11'b11111111111, 11'b11111110110, 11'b00000001010, 11'b00000000011, 11'b00000001111, 11'b00000000010, 11'b00000000001, 11'b11111110110, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b00000000110, 11'b00000000101, 11'b00000001001, 11'b11111111111, 11'b11111110110, 11'b00000000000, 11'b00000000000, 11'b00000001010, 11'b11111111001, 11'b11111101110, 11'b00000010001, 11'b11111110110, 11'b00000100101, 11'b11111111111, 11'b11111110100}, 
{11'b11111101101, 11'b11111111111, 11'b11111110010, 11'b00000000111, 11'b00000001000, 11'b11111111100, 11'b00000010000, 11'b11111111010, 11'b11111110000, 11'b11111110100, 11'b11111110111, 11'b11111110000, 11'b11111111000, 11'b00000000110, 11'b00000000000, 11'b00000000000, 11'b00000011010, 11'b11111111110, 11'b11111111111, 11'b00000001101, 11'b00000001001, 11'b11111101101, 11'b11111110011, 11'b00000000110, 11'b11111110010, 11'b11111111111, 11'b11111110111, 11'b11111110101, 11'b11111110010, 11'b00000001001, 11'b00000000111, 11'b11111111011, 11'b11111111101, 11'b11111100000, 11'b11111111010, 11'b00000000001, 11'b11111111011, 11'b11111110110, 11'b11111111111, 11'b00000000011, 11'b11111111100, 11'b11111111111, 11'b11111111110, 11'b11111101010, 11'b00000000000, 11'b00000000000, 11'b00000001010, 11'b11111111100, 11'b00000001101, 11'b11111111001, 11'b00000001001, 11'b11111111111, 11'b00000000111, 11'b11111110011, 11'b11111111111, 11'b00000010000, 11'b00000001010, 11'b00000001001, 11'b00000000000, 11'b11111110011, 11'b11111110110, 11'b11111101010, 11'b11111111111, 11'b00000000011}, 
{11'b00000001001, 11'b00000000000, 11'b00000000100, 11'b11111111111, 11'b00000000100, 11'b11111111011, 11'b00000000111, 11'b00000000001, 11'b00000000100, 11'b00000001010, 11'b11111110111, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b11111101010, 11'b11111110110, 11'b00000010100, 11'b11111111111, 11'b11111111110, 11'b00000000000, 11'b11111110011, 11'b00000000000, 11'b00000001000, 11'b00000000001, 11'b00000000001, 11'b00000001010, 11'b00000000000, 11'b00000000001, 11'b00000000000, 11'b11111111110, 11'b11111111001, 11'b11111101010, 11'b00000001000, 11'b00000001010, 11'b11111111111, 11'b11111111000, 11'b00000000000, 11'b11111101011, 11'b11111111110, 11'b11111111111, 11'b00000000110, 11'b11111111011, 11'b11111111111, 11'b00000011011, 11'b00000001110, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b11111111000, 11'b00000000100, 11'b00000000100, 11'b00000000101, 11'b00000000101, 11'b00000001100, 11'b00000001011, 11'b00000010101, 11'b11111111011, 11'b00000001100, 11'b00000000100, 11'b11111110101, 11'b00000000011, 11'b11111110011, 11'b11111110001, 11'b11111110000}, 
{11'b00000000000, 11'b00000000111, 11'b11111111001, 11'b00000000000, 11'b11111111110, 11'b11111111110, 11'b11111101010, 11'b11111111111, 11'b00000001000, 11'b00000000111, 11'b00000000111, 11'b11111110011, 11'b11111111101, 11'b00000001001, 11'b11111111111, 11'b00000000000, 11'b11111100101, 11'b11111111111, 11'b00000001011, 11'b00000000010, 11'b00000000111, 11'b11111111100, 11'b00000000111, 11'b00000001100, 11'b11111110100, 11'b11111110111, 11'b11111111111, 11'b11111111101, 11'b00000000010, 11'b00000000000, 11'b11111111111, 11'b00000001010, 11'b11111101000, 11'b00000001011, 11'b00000010000, 11'b00000000011, 11'b00000000011, 11'b11111111100, 11'b00000000011, 11'b11111111100, 11'b11111110111, 11'b11111111110, 11'b00000000101, 11'b00000010110, 11'b11111100100, 11'b11111110001, 11'b00000000110, 11'b11111111100, 11'b00000001110, 11'b11111111000, 11'b11111110101, 11'b11111110111, 11'b11111111111, 11'b00000000011, 11'b11111111010, 11'b11111100101, 11'b11111111011, 11'b11111111111, 11'b00000000001, 11'b11111101100, 11'b00000100011, 11'b11111101110, 11'b00000010001, 11'b00000000100}, 
{11'b00000000010, 11'b11111111001, 11'b00000010100, 11'b11111110110, 11'b11111110001, 11'b00000000010, 11'b00000001001, 11'b00000001001, 11'b11111111010, 11'b11111111010, 11'b00000000001, 11'b00000000111, 11'b00000000111, 11'b00000000001, 11'b11111111001, 11'b00000000100, 11'b00000001111, 11'b11111111111, 11'b11111110111, 11'b00000000000, 11'b00000000010, 11'b00000000000, 11'b11111110110, 11'b00000000011, 11'b00000011001, 11'b00000000000, 11'b00000000101, 11'b11111100110, 11'b11111111101, 11'b00000000000, 11'b11111111001, 11'b11111110110, 11'b00000001110, 11'b11111111111, 11'b11111111110, 11'b11111110110, 11'b00000000100, 11'b00000001001, 11'b11111111111, 11'b11111111110, 11'b11111111010, 11'b00000000111, 11'b00000000000, 11'b11111101010, 11'b00000001001, 11'b00000001100, 11'b11111111111, 11'b00000000000, 11'b11111110010, 11'b11111111101, 11'b11111111111, 11'b11111110101, 11'b00000000000, 11'b11111111010, 11'b00000000001, 11'b11111100101, 11'b11111111111, 11'b11111111111, 11'b00000001000, 11'b00000010010, 11'b11111101001, 11'b00000010000, 11'b00000000001, 11'b11111111101}, 
{11'b00000001001, 11'b00000100111, 11'b00000001111, 11'b00000001001, 11'b11111110000, 11'b11111110101, 11'b11110101100, 11'b11111110001, 11'b00000001100, 11'b11111111111, 11'b00000001001, 11'b00000011011, 11'b00000000010, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b11111111001, 11'b11111111001, 11'b00000000111, 11'b11111101111, 11'b11111101010, 11'b11111111100, 11'b11111101101, 11'b00000000000, 11'b11110110111, 11'b00000011010, 11'b00000011111, 11'b00000010011, 11'b11111001000, 11'b11111110101, 11'b11111101001, 11'b11111100101, 11'b11110101111, 11'b00000010101, 11'b11111111110, 11'b00000001010, 11'b00000000000, 11'b11111010010, 11'b00000000000, 11'b00000000000, 11'b00000000001, 11'b00000100000, 11'b11111111001, 11'b11111101011, 11'b00000011100, 11'b11111110001, 11'b11111110101, 11'b11111110011, 11'b00000001111, 11'b00000010001, 11'b11111111101, 11'b11111110100, 11'b11111111111, 11'b11111111100, 11'b00000000000, 11'b11111110011, 11'b00000010011, 11'b00000100010, 11'b00000010110, 11'b11111100010, 11'b11110001001, 11'b00000011100, 11'b00000000010, 11'b00000001010}, 
{11'b11111111000, 11'b00000001010, 11'b00000001010, 11'b11111111111, 11'b11111110100, 11'b11111111101, 11'b11111110011, 11'b11111111110, 11'b00000000100, 11'b11111111101, 11'b11111111111, 11'b11111111110, 11'b11111111111, 11'b11111111010, 11'b11111111111, 11'b11111111100, 11'b00000001010, 11'b11111111111, 11'b11111101011, 11'b00000001110, 11'b00000010011, 11'b00000001101, 11'b11111110101, 11'b11111111011, 11'b11111110100, 11'b11111110110, 11'b00000000111, 11'b00000000111, 11'b00000000111, 11'b00000001011, 11'b00000000001, 11'b00000001100, 11'b11111111110, 11'b00000000000, 11'b00000001001, 11'b00000000100, 11'b11111111101, 11'b11111111111, 11'b00000000000, 11'b11111110110, 11'b11111111000, 11'b11111111100, 11'b11111110100, 11'b00000001110, 11'b00000000000, 11'b11111111111, 11'b11111111101, 11'b11111111011, 11'b11111100110, 11'b11111111110, 11'b11111111000, 11'b11111111011, 11'b11111111100, 11'b00000001000, 11'b00000010101, 11'b00000000101, 11'b11111111111, 11'b11111110101, 11'b11111111111, 11'b00000000000, 11'b00000001010, 11'b11111111111, 11'b00000000001, 11'b00000000000}
};

localparam logic signed [10:0] bias [64] = '{
11'b11111111110,  // -0.037350185215473175
11'b00000001000,  // 0.27355897426605225
11'b11111111100,  // -0.12378914654254913
11'b11111111101,  // -0.064457006752491
11'b00000000001,  // 0.05452875792980194
11'b00000000011,  // 0.11671770364046097
11'b00000000100,  // 0.13640816509723663
11'b00000000010,  // 0.07482525706291199
11'b00000000001,  // 0.04674031585454941
11'b11111111001,  // -0.20146161317825317
11'b11111111100,  // -0.09910125285387039
11'b00000000100,  // 0.15104414522647858
11'b11111111100,  // -0.10221704095602036
11'b11111111011,  // -0.1461549550294876
11'b11111111101,  // -0.08641516417264938
11'b00000000101,  // 0.16613510251045227
11'b11111111101,  // -0.0836295336484909
11'b11111111110,  // -0.05756539851427078
11'b11111111110,  // -0.03229188174009323
11'b11111111111,  // -0.028388574719429016
11'b00000000100,  // 0.1260243058204651
11'b11111111110,  // -0.037064336240291595
11'b00000000110,  // 0.19336333870887756
11'b00000000000,  // 0.02124214917421341
11'b00000001111,  // 0.4985624849796295
11'b00000000000,  // 0.0158411655575037
11'b11111111101,  // -0.08296407759189606
11'b00000000011,  // 0.11056788265705109
11'b00000000000,  // 0.01173810102045536
11'b11111111100,  // -0.10843746364116669
11'b00000001000,  // 0.27439257502555847
11'b00000000010,  // 0.09199801832437515
11'b00000001000,  // 0.27419957518577576
11'b00000001000,  // 0.27063727378845215
11'b11111111000,  // -0.24828937649726868
11'b00000000010,  // 0.07818280160427094
11'b11111111111,  // -0.005749030504375696
11'b00000000011,  // 0.10850494354963303
11'b00000000100,  // 0.13591453433036804
11'b11111111100,  // -0.12088628858327866
11'b11111111110,  // -0.05666546896100044
11'b00000000010,  // 0.09311636537313461
11'b00000000001,  // 0.05477767437696457
11'b00000000000,  // 0.029585206881165504
11'b11111110110,  // -0.31209176778793335
11'b11111111101,  // -0.08465463668107986
11'b11111111010,  // -0.16775836050510406
11'b00000000100,  // 0.14762157201766968
11'b11111111000,  // -0.23618532717227936
11'b00000000010,  // 0.06535740196704865
11'b11111111011,  // -0.12853026390075684
11'b11111111011,  // -0.13802281022071838
11'b11111111011,  // -0.15156887471675873
11'b00000000010,  // 0.07979883998632431
11'b00000000101,  // 0.18141601979732513
11'b11111111110,  // -0.054039113223552704
11'b11111111111,  // -0.010052933357656002
11'b00000000010,  // 0.06611225008964539
11'b00000000001,  // 0.05053366720676422
11'b00000000000,  // 0.026860840618610382
11'b00000000001,  // 0.03283466026186943
11'b00000000100,  // 0.15558314323425293
11'b11111110110,  // -0.2863388657569885
11'b11111111101   // -0.08769102394580841
};
endpackage