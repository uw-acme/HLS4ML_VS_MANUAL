// Width: 12
// NFRAC: 6
package dense_1_12_6;

localparam logic signed [11:0] weights [16][64] = '{ 
{12'b000000010000, 12'b111111010110, 12'b111111110100, 12'b111111110001, 12'b111111100110, 12'b000000000111, 12'b111110111101, 12'b000000000000, 12'b000000000011, 12'b000000010000, 12'b000000000000, 12'b111111100110, 12'b111111111111, 12'b000000001101, 12'b000000000010, 12'b111111101111, 12'b000000001110, 12'b000000000011, 12'b000000000000, 12'b111111111111, 12'b000000011000, 12'b111111101010, 12'b111111111110, 12'b000000011110, 12'b111111101011, 12'b111111010100, 12'b111111101110, 12'b111111110011, 12'b111111111001, 12'b111111111111, 12'b000000000010, 12'b000000001111, 12'b000000001100, 12'b111111111111, 12'b000000000000, 12'b000000010011, 12'b111111111110, 12'b111111101111, 12'b000000000001, 12'b000000001100, 12'b111111111111, 12'b000000010001, 12'b111111101110, 12'b000000111011, 12'b111111111111, 12'b000000011100, 12'b000000000000, 12'b000000001011, 12'b000000001100, 12'b111111111110, 12'b000000000000, 12'b000000001010, 12'b000000001101, 12'b000000000100, 12'b111111111000, 12'b111111101100, 12'b000000100010, 12'b111111100000, 12'b000000011101, 12'b111111101001, 12'b000000110010, 12'b111111111111, 12'b000000000000, 12'b000000000101}, 
{12'b000000000000, 12'b111111101011, 12'b111111110111, 12'b111111101110, 12'b111111101011, 12'b000000000110, 12'b111111001111, 12'b111111111111, 12'b111111110001, 12'b000000001011, 12'b000000000000, 12'b111111111010, 12'b000000001100, 12'b000000000000, 12'b111111111111, 12'b000000001101, 12'b111111111111, 12'b000000000000, 12'b111111110100, 12'b111111101111, 12'b000000011100, 12'b111111111010, 12'b000000000011, 12'b000000101100, 12'b000000010000, 12'b111111110001, 12'b111111110001, 12'b111111111111, 12'b111111111001, 12'b111111100110, 12'b111111111100, 12'b000000011101, 12'b000000010001, 12'b000000100011, 12'b000000101000, 12'b000000000011, 12'b111111111000, 12'b111111100100, 12'b000000000011, 12'b000000001100, 12'b000000000001, 12'b000000001101, 12'b111111110010, 12'b000000010000, 12'b000000001011, 12'b000000000011, 12'b111111101010, 12'b000000000101, 12'b000000010000, 12'b000000000001, 12'b000000000001, 12'b000001001010, 12'b111111111011, 12'b111111111001, 12'b111111111100, 12'b111111111111, 12'b000000010000, 12'b111111101000, 12'b000000111111, 12'b000000000000, 12'b000000100001, 12'b000000001111, 12'b000000110100, 12'b000000001001}, 
{12'b111111111111, 12'b000000000000, 12'b111111111010, 12'b111111110100, 12'b111111110100, 12'b000000000010, 12'b000001011110, 12'b111111111111, 12'b111110101110, 12'b111111111111, 12'b111111111111, 12'b111111111110, 12'b111111110001, 12'b000000000000, 12'b111111111111, 12'b000000001010, 12'b000000111001, 12'b111111111111, 12'b000000000100, 12'b000000000000, 12'b000000011010, 12'b111111010001, 12'b000000100100, 12'b111111010010, 12'b000000111100, 12'b111111101001, 12'b111111110000, 12'b111111010010, 12'b000001010001, 12'b000000010001, 12'b000000000000, 12'b000000100001, 12'b000001000001, 12'b111110110011, 12'b111111111001, 12'b000000000010, 12'b111111110001, 12'b000000111001, 12'b111111111101, 12'b000000010100, 12'b000000010101, 12'b000000010111, 12'b111111111111, 12'b111111111111, 12'b111111111110, 12'b000000001010, 12'b111111101110, 12'b111111110101, 12'b111111111110, 12'b000000011001, 12'b111111110100, 12'b000000001001, 12'b111111111111, 12'b000000001000, 12'b111111110100, 12'b111111111111, 12'b111111101100, 12'b111111010101, 12'b111111111111, 12'b000000000000, 12'b000001100010, 12'b000000000000, 12'b111111111111, 12'b111111101100}, 
{12'b111111100010, 12'b111111101000, 12'b111111010011, 12'b000000010011, 12'b111111101011, 12'b111110101001, 12'b111111111000, 12'b111111101100, 12'b000000001110, 12'b111111111111, 12'b000001010000, 12'b111111111001, 12'b111111001101, 12'b000000100101, 12'b000000000001, 12'b111111111111, 12'b111111100011, 12'b111111111111, 12'b000000000000, 12'b111111110001, 12'b111110110110, 12'b111111111000, 12'b111111010011, 12'b000000001100, 12'b111111100111, 12'b111111000101, 12'b000000010100, 12'b000000101111, 12'b000001010010, 12'b111111100010, 12'b111111011010, 12'b000000000100, 12'b000000100000, 12'b111111001010, 12'b111111101011, 12'b000000000000, 12'b111111010001, 12'b000000001111, 12'b111111100011, 12'b000000000111, 12'b000000011101, 12'b000000001010, 12'b000000000000, 12'b000000000001, 12'b000000100011, 12'b111111110011, 12'b111111111111, 12'b111111101001, 12'b111111111111, 12'b111111111001, 12'b111111011000, 12'b000000000101, 12'b111111111111, 12'b000000001101, 12'b000000010100, 12'b000000101001, 12'b111111000010, 12'b111111000100, 12'b111111010010, 12'b000000110111, 12'b000001101111, 12'b111111000110, 12'b111111111100, 12'b000000011011}, 
{12'b000000010101, 12'b111111011000, 12'b111111101111, 12'b111111111111, 12'b111111110110, 12'b000000010101, 12'b000000001100, 12'b111111111111, 12'b111111011001, 12'b111111110000, 12'b111111101000, 12'b000000000011, 12'b000000000000, 12'b000000000000, 12'b111111111101, 12'b000000010110, 12'b000000001000, 12'b111111100110, 12'b000000000001, 12'b000000000000, 12'b000000001101, 12'b111111111000, 12'b000000000100, 12'b111111111110, 12'b000001000100, 12'b111111110100, 12'b111111101110, 12'b111111100110, 12'b000000000000, 12'b000000001010, 12'b000000000111, 12'b000000010001, 12'b111111111111, 12'b000000000100, 12'b000000001000, 12'b111111111111, 12'b000000000000, 12'b000000111000, 12'b111111101101, 12'b111111111011, 12'b000000011011, 12'b000000001111, 12'b111111100000, 12'b000000000000, 12'b111110111011, 12'b111111111111, 12'b111111111000, 12'b000000000000, 12'b111111111111, 12'b111111111110, 12'b111111111111, 12'b000000001100, 12'b111111111111, 12'b000000010100, 12'b111111110011, 12'b111111010000, 12'b111111100010, 12'b111111011111, 12'b111111011000, 12'b000000101111, 12'b000001010111, 12'b000000110010, 12'b000000000111, 12'b111111111111}, 
{12'b111111100011, 12'b111111010111, 12'b000000000000, 12'b000000010011, 12'b000000010010, 12'b111111110010, 12'b000000100101, 12'b111111111111, 12'b000000001111, 12'b111111111111, 12'b111111111111, 12'b111111111011, 12'b111111110100, 12'b000000100101, 12'b111111111010, 12'b000000000000, 12'b111111011000, 12'b111111101001, 12'b000000000000, 12'b111111111111, 12'b111111111100, 12'b111111101011, 12'b111111101011, 12'b000000011101, 12'b111111101011, 12'b111111111111, 12'b000000010000, 12'b111111111011, 12'b111111000100, 12'b111111111111, 12'b111111111011, 12'b111111111111, 12'b111111111111, 12'b000000000010, 12'b000000001000, 12'b000000010110, 12'b000000000000, 12'b111111111001, 12'b111111101111, 12'b111111111111, 12'b111111110101, 12'b111111011110, 12'b000000011001, 12'b000000000000, 12'b000000100110, 12'b000000000000, 12'b111111111111, 12'b000000000110, 12'b111111100101, 12'b000000001110, 12'b000000000000, 12'b111111111001, 12'b111111101000, 12'b000000011000, 12'b111111111111, 12'b000000010110, 12'b000000001101, 12'b000000001101, 12'b111111111110, 12'b111111111111, 12'b111111001100, 12'b111111110111, 12'b111111111100, 12'b111111111111}, 
{12'b111111101101, 12'b111111101010, 12'b111111100100, 12'b111111111011, 12'b111111110111, 12'b000000000110, 12'b111111010011, 12'b111111110110, 12'b111111110001, 12'b111111111111, 12'b111111101101, 12'b000000010110, 12'b000000000010, 12'b000000001000, 12'b000000010011, 12'b000000000000, 12'b000000110011, 12'b000000000101, 12'b000000001111, 12'b000000010001, 12'b111111110101, 12'b000000010111, 12'b111111110000, 12'b111111011111, 12'b000000001011, 12'b000000100001, 12'b111111111111, 12'b000000000011, 12'b111111000011, 12'b000000010010, 12'b000000010001, 12'b111111101000, 12'b000000011110, 12'b000000101010, 12'b000000000000, 12'b000000010101, 12'b111111111111, 12'b000000010010, 12'b000000001100, 12'b000000000000, 12'b111111111000, 12'b111111101000, 12'b000000001001, 12'b000000011110, 12'b000000100001, 12'b111111110101, 12'b111111111010, 12'b111111110011, 12'b111111110111, 12'b000000000111, 12'b000000000000, 12'b000000000010, 12'b000000000000, 12'b000000001011, 12'b111111110100, 12'b000000110001, 12'b000000010110, 12'b111111111110, 12'b000000011000, 12'b000000001101, 12'b111110010111, 12'b111111011011, 12'b111111110100, 12'b111111111111}, 
{12'b000000000000, 12'b000000001111, 12'b111111111111, 12'b111111111111, 12'b111111101011, 12'b111111111110, 12'b111111101111, 12'b000000000000, 12'b000000000001, 12'b000000011000, 12'b000000000000, 12'b111111100111, 12'b111111111011, 12'b000000000000, 12'b111111111100, 12'b111111100011, 12'b111111001001, 12'b111111111111, 12'b111111011001, 12'b111111100011, 12'b111111100111, 12'b000000010110, 12'b000000000011, 12'b111111110110, 12'b111111100100, 12'b000000001001, 12'b000000000000, 12'b000000011111, 12'b000000110011, 12'b111111111101, 12'b000000000000, 12'b000000001110, 12'b111111010100, 12'b111111101000, 12'b000000000011, 12'b000000000101, 12'b111111101110, 12'b000000001111, 12'b000000001000, 12'b111111110110, 12'b111111100101, 12'b111111111101, 12'b000000000010, 12'b111111110101, 12'b000000000011, 12'b000000001110, 12'b111111111000, 12'b000000000001, 12'b000000000000, 12'b111111110010, 12'b111111100111, 12'b000000011010, 12'b000000001000, 12'b111111110100, 12'b000000001000, 12'b111111111100, 12'b111111100001, 12'b111111110111, 12'b111111111100, 12'b111111111011, 12'b000000110101, 12'b000000001100, 12'b111111111100, 12'b111111111111}, 
{12'b000000000000, 12'b000000100101, 12'b111111011010, 12'b111111110001, 12'b000000010100, 12'b111111110010, 12'b000001001101, 12'b111111101101, 12'b111111111111, 12'b000000010010, 12'b000000010000, 12'b111111111111, 12'b111111111100, 12'b111111100001, 12'b000000010010, 12'b000000001010, 12'b111111110011, 12'b111111111111, 12'b000000000000, 12'b000000000000, 12'b000000010000, 12'b111111100010, 12'b000000011001, 12'b000000100111, 12'b111111111010, 12'b111111111111, 12'b111111111110, 12'b111111111111, 12'b000000101111, 12'b000000000000, 12'b111111101110, 12'b000000000000, 12'b000000011000, 12'b111111001100, 12'b111111011101, 12'b000000001100, 12'b000000001000, 12'b111111011011, 12'b111111110011, 12'b111111110010, 12'b000000011001, 12'b000000011001, 12'b000000000000, 12'b111111101110, 12'b000000000000, 12'b000000011001, 12'b111111111100, 12'b111111111111, 12'b000000000000, 12'b000000001111, 12'b111111111100, 12'b111111110011, 12'b000000010110, 12'b111111110010, 12'b000000010001, 12'b000000100101, 12'b000000000010, 12'b000000010000, 12'b111111100110, 12'b111111101000, 12'b000000110101, 12'b111111110111, 12'b000000000010, 12'b111111111010}, 
{12'b000000000001, 12'b111111100011, 12'b000000010111, 12'b111111101101, 12'b111111111111, 12'b000000001101, 12'b111111011010, 12'b000000001100, 12'b000000011111, 12'b000000001001, 12'b000000010111, 12'b000000010100, 12'b111111101100, 12'b111111111011, 12'b111111111100, 12'b000000000000, 12'b111111000010, 12'b000000010100, 12'b111111111101, 12'b000000000001, 12'b111111101001, 12'b000000000100, 12'b000000001001, 12'b111111111111, 12'b111111100010, 12'b111111111100, 12'b111111111010, 12'b000001001111, 12'b111111010101, 12'b000000000100, 12'b000000000110, 12'b111111111100, 12'b111111110001, 12'b000000000111, 12'b111111111010, 12'b111111110111, 12'b111111110100, 12'b111111110010, 12'b111111111110, 12'b111111101100, 12'b000000010100, 12'b000000000111, 12'b000000011111, 12'b000000000101, 12'b000000000010, 12'b111111101101, 12'b000000000000, 12'b111111111111, 12'b111111111111, 12'b000000001100, 12'b000000001011, 12'b000000010010, 12'b111111111111, 12'b111111101101, 12'b000000000000, 12'b000000000000, 12'b000000010100, 12'b111111110011, 12'b111111011100, 12'b000000100011, 12'b111111101101, 12'b000001001010, 12'b111111111110, 12'b111111101001}, 
{12'b111111011011, 12'b111111111111, 12'b111111100101, 12'b000000001110, 12'b000000010000, 12'b111111111001, 12'b000000100001, 12'b111111110101, 12'b111111100001, 12'b111111101000, 12'b111111101111, 12'b111111100001, 12'b111111110001, 12'b000000001100, 12'b000000000000, 12'b000000000000, 12'b000000110101, 12'b111111111101, 12'b111111111111, 12'b000000011010, 12'b000000010010, 12'b111111011010, 12'b111111100111, 12'b000000001100, 12'b111111100100, 12'b111111111110, 12'b111111101111, 12'b111111101010, 12'b111111100100, 12'b000000010011, 12'b000000001110, 12'b111111110110, 12'b111111111011, 12'b111111000001, 12'b111111110100, 12'b000000000011, 12'b111111110111, 12'b111111101101, 12'b111111111111, 12'b000000000111, 12'b111111111000, 12'b111111111111, 12'b111111111101, 12'b111111010101, 12'b000000000000, 12'b000000000000, 12'b000000010101, 12'b111111111000, 12'b000000011011, 12'b111111110011, 12'b000000010010, 12'b111111111111, 12'b000000001110, 12'b111111100110, 12'b111111111111, 12'b000000100000, 12'b000000010100, 12'b000000010010, 12'b000000000001, 12'b111111100110, 12'b111111101100, 12'b111111010100, 12'b111111111111, 12'b000000000110}, 
{12'b000000010011, 12'b000000000000, 12'b000000001000, 12'b111111111111, 12'b000000001001, 12'b111111110111, 12'b000000001111, 12'b000000000010, 12'b000000001000, 12'b000000010101, 12'b111111101111, 12'b111111111110, 12'b111111111111, 12'b111111111111, 12'b111111010101, 12'b111111101100, 12'b000000101000, 12'b111111111110, 12'b111111111100, 12'b000000000000, 12'b111111100111, 12'b000000000000, 12'b000000010000, 12'b000000000010, 12'b000000000010, 12'b000000010101, 12'b000000000000, 12'b000000000010, 12'b000000000000, 12'b111111111100, 12'b111111110011, 12'b111111010101, 12'b000000010000, 12'b000000010101, 12'b111111111110, 12'b111111110000, 12'b000000000000, 12'b111111010110, 12'b111111111101, 12'b111111111111, 12'b000000001100, 12'b111111110111, 12'b111111111111, 12'b000000110110, 12'b000000011100, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111110000, 12'b000000001001, 12'b000000001001, 12'b000000001011, 12'b000000001010, 12'b000000011000, 12'b000000010110, 12'b000000101010, 12'b111111110111, 12'b000000011001, 12'b000000001001, 12'b111111101011, 12'b000000000111, 12'b111111100111, 12'b111111100011, 12'b111111100000}, 
{12'b000000000000, 12'b000000001110, 12'b111111110011, 12'b000000000000, 12'b111111111100, 12'b111111111101, 12'b111111010101, 12'b111111111111, 12'b000000010000, 12'b000000001111, 12'b000000001111, 12'b111111100110, 12'b111111111010, 12'b000000010010, 12'b111111111111, 12'b000000000000, 12'b111111001010, 12'b111111111111, 12'b000000010111, 12'b000000000100, 12'b000000001111, 12'b111111111000, 12'b000000001111, 12'b000000011001, 12'b111111101001, 12'b111111101110, 12'b111111111111, 12'b111111111010, 12'b000000000100, 12'b000000000000, 12'b111111111111, 12'b000000010100, 12'b111111010000, 12'b000000010111, 12'b000000100000, 12'b000000000111, 12'b000000000111, 12'b111111111001, 12'b000000000111, 12'b111111111001, 12'b111111101111, 12'b111111111100, 12'b000000001010, 12'b000000101100, 12'b111111001001, 12'b111111100011, 12'b000000001100, 12'b111111111001, 12'b000000011100, 12'b111111110000, 12'b111111101010, 12'b111111101110, 12'b111111111111, 12'b000000000111, 12'b111111110101, 12'b111111001010, 12'b111111110110, 12'b111111111111, 12'b000000000010, 12'b111111011000, 12'b000001000111, 12'b111111011101, 12'b000000100010, 12'b000000001001}, 
{12'b000000000101, 12'b111111110011, 12'b000000101000, 12'b111111101100, 12'b111111100010, 12'b000000000101, 12'b000000010011, 12'b000000010011, 12'b111111110100, 12'b111111110101, 12'b000000000011, 12'b000000001110, 12'b000000001111, 12'b000000000011, 12'b111111110010, 12'b000000001000, 12'b000000011110, 12'b111111111111, 12'b111111101110, 12'b000000000000, 12'b000000000100, 12'b000000000001, 12'b111111101101, 12'b000000000111, 12'b000000110010, 12'b000000000000, 12'b000000001011, 12'b111111001101, 12'b111111111011, 12'b000000000000, 12'b111111110011, 12'b111111101100, 12'b000000011101, 12'b111111111110, 12'b111111111101, 12'b111111101100, 12'b000000001000, 12'b000000010010, 12'b111111111111, 12'b111111111101, 12'b111111110100, 12'b000000001110, 12'b000000000000, 12'b111111010100, 12'b000000010011, 12'b000000011001, 12'b111111111111, 12'b000000000001, 12'b111111100100, 12'b111111111011, 12'b111111111111, 12'b111111101011, 12'b000000000000, 12'b111111110100, 12'b000000000011, 12'b111111001011, 12'b111111111111, 12'b111111111111, 12'b000000010001, 12'b000000100100, 12'b111111010011, 12'b000000100001, 12'b000000000010, 12'b111111111011}, 
{12'b000000010010, 12'b000001001111, 12'b000000011111, 12'b000000010010, 12'b111111100001, 12'b111111101011, 12'b111101011001, 12'b111111100010, 12'b000000011001, 12'b111111111111, 12'b000000010010, 12'b000000110111, 12'b000000000100, 12'b000000000000, 12'b111111111110, 12'b000000000000, 12'b111111110011, 12'b111111110011, 12'b000000001110, 12'b111111011111, 12'b111111010101, 12'b111111111001, 12'b111111011010, 12'b000000000001, 12'b111101101110, 12'b000000110100, 12'b000000111111, 12'b000000100110, 12'b111110010000, 12'b111111101011, 12'b111111010011, 12'b111111001010, 12'b111101011110, 12'b000000101011, 12'b111111111101, 12'b000000010100, 12'b000000000001, 12'b111110100100, 12'b000000000000, 12'b000000000000, 12'b000000000010, 12'b000001000001, 12'b111111110010, 12'b111111010110, 12'b000000111001, 12'b111111100011, 12'b111111101011, 12'b111111100110, 12'b000000011110, 12'b000000100010, 12'b111111111011, 12'b111111101001, 12'b111111111111, 12'b111111111000, 12'b000000000000, 12'b111111100111, 12'b000000100110, 12'b000001000101, 12'b000000101101, 12'b111111000101, 12'b111100010011, 12'b000000111000, 12'b000000000101, 12'b000000010100}, 
{12'b111111110000, 12'b000000010101, 12'b000000010100, 12'b111111111111, 12'b111111101000, 12'b111111111010, 12'b111111100111, 12'b111111111100, 12'b000000001001, 12'b111111111011, 12'b111111111110, 12'b111111111101, 12'b111111111111, 12'b111111110100, 12'b111111111110, 12'b111111111001, 12'b000000010100, 12'b111111111111, 12'b111111010110, 12'b000000011101, 12'b000000100110, 12'b000000011010, 12'b111111101011, 12'b111111110111, 12'b111111101001, 12'b111111101101, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000010111, 12'b000000000010, 12'b000000011000, 12'b111111111101, 12'b000000000000, 12'b000000010011, 12'b000000001000, 12'b111111111011, 12'b111111111111, 12'b000000000000, 12'b111111101101, 12'b111111110001, 12'b111111111000, 12'b111111101001, 12'b000000011100, 12'b000000000000, 12'b111111111111, 12'b111111111010, 12'b111111110110, 12'b111111001100, 12'b111111111101, 12'b111111110001, 12'b111111110110, 12'b111111111001, 12'b000000010000, 12'b000000101011, 12'b000000001011, 12'b111111111111, 12'b111111101010, 12'b111111111110, 12'b000000000000, 12'b000000010100, 12'b111111111110, 12'b000000000010, 12'b000000000000}
};

localparam logic signed [11:0] bias [64] = '{
12'b111111111101,  // -0.037350185215473175
12'b000000010001,  // 0.27355897426605225
12'b111111111000,  // -0.12378914654254913
12'b111111111011,  // -0.064457006752491
12'b000000000011,  // 0.05452875792980194
12'b000000000111,  // 0.11671770364046097
12'b000000001000,  // 0.13640816509723663
12'b000000000100,  // 0.07482525706291199
12'b000000000010,  // 0.04674031585454941
12'b111111110011,  // -0.20146161317825317
12'b111111111001,  // -0.09910125285387039
12'b000000001001,  // 0.15104414522647858
12'b111111111001,  // -0.10221704095602036
12'b111111110110,  // -0.1461549550294876
12'b111111111010,  // -0.08641516417264938
12'b000000001010,  // 0.16613510251045227
12'b111111111010,  // -0.0836295336484909
12'b111111111100,  // -0.05756539851427078
12'b111111111101,  // -0.03229188174009323
12'b111111111110,  // -0.028388574719429016
12'b000000001000,  // 0.1260243058204651
12'b111111111101,  // -0.037064336240291595
12'b000000001100,  // 0.19336333870887756
12'b000000000001,  // 0.02124214917421341
12'b000000011111,  // 0.4985624849796295
12'b000000000001,  // 0.0158411655575037
12'b111111111010,  // -0.08296407759189606
12'b000000000111,  // 0.11056788265705109
12'b000000000000,  // 0.01173810102045536
12'b111111111001,  // -0.10843746364116669
12'b000000010001,  // 0.27439257502555847
12'b000000000101,  // 0.09199801832437515
12'b000000010001,  // 0.27419957518577576
12'b000000010001,  // 0.27063727378845215
12'b111111110000,  // -0.24828937649726868
12'b000000000101,  // 0.07818280160427094
12'b111111111111,  // -0.005749030504375696
12'b000000000110,  // 0.10850494354963303
12'b000000001000,  // 0.13591453433036804
12'b111111111000,  // -0.12088628858327866
12'b111111111100,  // -0.05666546896100044
12'b000000000101,  // 0.09311636537313461
12'b000000000011,  // 0.05477767437696457
12'b000000000001,  // 0.029585206881165504
12'b111111101100,  // -0.31209176778793335
12'b111111111010,  // -0.08465463668107986
12'b111111110101,  // -0.16775836050510406
12'b000000001001,  // 0.14762157201766968
12'b111111110000,  // -0.23618532717227936
12'b000000000100,  // 0.06535740196704865
12'b111111110111,  // -0.12853026390075684
12'b111111110111,  // -0.13802281022071838
12'b111111110110,  // -0.15156887471675873
12'b000000000101,  // 0.07979883998632431
12'b000000001011,  // 0.18141601979732513
12'b111111111100,  // -0.054039113223552704
12'b111111111111,  // -0.010052933357656002
12'b000000000100,  // 0.06611225008964539
12'b000000000011,  // 0.05053366720676422
12'b000000000001,  // 0.026860840618610382
12'b000000000010,  // 0.03283466026186943
12'b000000001001,  // 0.15558314323425293
12'b111111101101,  // -0.2863388657569885
12'b111111111010   // -0.08769102394580841
};
endpackage