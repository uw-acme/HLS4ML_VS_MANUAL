//Width: 25
//Int: 9
package dense_3_gen;

localparam logic signed [24:0] weights [32][32] = '{
{25'b1111111111111001101101101, 25'b1111111111001000000010010, 25'b1111111111001100000100111, 25'b1111111111100111100111111, 25'b0000000000101011111011011, 25'b0000000000000101100111101, 25'b1111111111111110010111001, 25'b1111111111111111111001011, 25'b1111111111111111111111110, 25'b1111111111111111111110100, 25'b0000000000010000001000111, 25'b1111111110111100100011111, 25'b1111111111111000010111000, 25'b0000000001101100011011011, 25'b1111111111100001000101101, 25'b1111111110001000100111011, 25'b1111111111111011010110001, 25'b0000000000001110010000111, 25'b0000000000110111101011010, 25'b1111111111010011011010111, 25'b1111111101110111100110001, 25'b1111111111111010000111111, 25'b0000000000000110010011011, 25'b1111111111001100011000010, 25'b0000000000000000000001101, 25'b0000000010000001100111100, 25'b1111111101000101100100110, 25'b1111111111100011101000010, 25'b1111111111001110010001010, 25'b1111111111101100110010100, 25'b0000000000110110001001110, 25'b1111111111101011100110101},
{25'b0000000001011111101101000, 25'b0000000011011101011100011, 25'b0000000000110011011101110, 25'b1111111110101011110100010, 25'b0000000000011111010001011, 25'b1111111111011101000000101, 25'b1111111111110010000111100, 25'b0000000010001011100000011, 25'b0000000000000000110001000, 25'b1111111111111111111111001, 25'b1111111111111011111100000, 25'b1111111110110100101101100, 25'b1111111111100110001110011, 25'b0000000001000101001010111, 25'b1111111011110010011101100, 25'b1111111111000011101011100, 25'b1111111111111111111111101, 25'b1111111111111110111100001, 25'b1111111111111001010000110, 25'b1111111111101010111110001, 25'b1111111111011110111011011, 25'b1111111111011100110000011, 25'b0000000000000010001101011, 25'b1111111111111111110010101, 25'b1111111111111111001011011, 25'b1111111101110110110001010, 25'b0000000000000001100000001, 25'b0000000000111100010010001, 25'b1111111111110111111001101, 25'b1111111110100111101101011, 25'b0000000000000000010110001, 25'b0000000000000100110110001},
{25'b1111111110000001111001001, 25'b0000000000010111100101000, 25'b0000000000000001010111111, 25'b0000000000101001010011100, 25'b1111111110101111010100011, 25'b0000000000000000000100001, 25'b0000000000000000001101100, 25'b1111111110010100100101110, 25'b0000000001000100100110010, 25'b1111111111011110011101110, 25'b1111111111011110110010101, 25'b1111111101000001101011100, 25'b1111111111011000001100111, 25'b0000000001000001011001100, 25'b0000000000100001110001010, 25'b1111111111111111110010010, 25'b1111111111110001010111010, 25'b1111111111111100111110011, 25'b1111111110010111101111011, 25'b0000000000000000011001101, 25'b0000000000001111111101010, 25'b0000000000001000110101001, 25'b0000000000011010110001110, 25'b0000000001110000101001101, 25'b0000000000000100110110000, 25'b1111111110011011000111110, 25'b0000000001100010001110001, 25'b0000000000000000000101101, 25'b0000000000010101001110101, 25'b1111111111111101001011110, 25'b0000000000000000000111110, 25'b0000000100100010011010101},
{25'b0000000001101011001110011, 25'b1111111111111111111111100, 25'b1111111111100111000111111, 25'b0000000010100111100000111, 25'b0000000010011101001100100, 25'b0000000000000000000010110, 25'b0000000000001001011011101, 25'b0000000001101000001010111, 25'b1111111111001101010100111, 25'b1111111111111111111110100, 25'b1111111110010110100111111, 25'b0000000000001111010100011, 25'b0000000000100010000111011, 25'b1111111110100000010101001, 25'b0000000000001011111110010, 25'b1111111111101011100010111, 25'b1111111111111111111111000, 25'b1111111111010001011001110, 25'b0000000000000100111011001, 25'b0000000000000111000100001, 25'b0000000000000010000010001, 25'b1111111111110110101010010, 25'b0000000010011000110010110, 25'b0000000001010111110001110, 25'b0000000001010100010100000, 25'b0000000000111111100010010, 25'b0000000001010111011100101, 25'b0000000000000000000011101, 25'b1111111111110000111001011, 25'b0000000001110011111111010, 25'b0000000000111111111000101, 25'b1111111111101001100001101},
{25'b0000000010000000000100000, 25'b1111111111110100000010110, 25'b1111111110100111010001110, 25'b1111111100111111100111000, 25'b0000000001111010001110100, 25'b0000000000000000000010001, 25'b1111111110010111000000000, 25'b1111111110110111101001101, 25'b1111111111110100000101001, 25'b1111111100110000110110000, 25'b1111111011100101001010110, 25'b0000000001111001000000110, 25'b0000000010101011001101010, 25'b0000000010000101111110010, 25'b1111111101101100110010110, 25'b1111111100111001100110100, 25'b0000000000000000000001000, 25'b1111111111011011110011001, 25'b0000000000110011011000110, 25'b0000000000100011100000101, 25'b1111111111001111110001110, 25'b1111111111111110010111111, 25'b0000000010111000110000000, 25'b1111111010100000000100010, 25'b0000000000010110100010001, 25'b1111111101010111011010000, 25'b0000000000010000110001110, 25'b1111111111000000011110101, 25'b1111111110110011100110100, 25'b1111111111111111111010111, 25'b0000000000010001111010110, 25'b0000000010010100100111100},
{25'b0000000000001011000011101, 25'b1111111111110101011010110, 25'b1111111110110001011001110, 25'b1111111110111101010111011, 25'b0000000001011111001010010, 25'b0000000000000000000010110, 25'b1111111110111000011000011, 25'b1111111111011101001001111, 25'b1111111110010010011001001, 25'b1111111111101111100110100, 25'b1111111111111111111000100, 25'b0000000000101001000010101, 25'b0000000000000000000000010, 25'b0000000001011011100101111, 25'b1111111101111110100001011, 25'b1111111111011111010100101, 25'b0000000000010110110011000, 25'b1111111110110100111111101, 25'b1111111111001101011011110, 25'b1111111111111111111110111, 25'b0000000000000011000111101, 25'b0000000001001100101110000, 25'b0000000001110111100011110, 25'b1111111111111101010001000, 25'b1111111111111111111001000, 25'b0000000001100110100101011, 25'b1111111101110011010101000, 25'b1111111111111111111110001, 25'b1111111111000011011100111, 25'b1111111111110110100100101, 25'b1111111111111111001100001, 25'b0000000000000001101010001},
{25'b0000000000010000101010001, 25'b1111111110101010111001111, 25'b0000000000011011101111100, 25'b1111111111110110001001110, 25'b1111111111111110000100101, 25'b0000000000100110110000110, 25'b1111111111100100110111111, 25'b1111111101010010101010110, 25'b1111111111111111111110100, 25'b1111111111001010101010100, 25'b1111111110001011000100111, 25'b0000000001111000111001000, 25'b0000000000000001110101000, 25'b0000000010101111001100111, 25'b0000000011010100001001010, 25'b0000000000000000101010101, 25'b1111111111111111111111110, 25'b1111111110101111010010000, 25'b1111111111110000001001011, 25'b0000000001000101111110111, 25'b1111111100111111111111000, 25'b0000000000100111111011101, 25'b0000000001010011100010001, 25'b0000000000000100110111100, 25'b0000000000100110011011111, 25'b0000000100111110010010001, 25'b1111111110011011000110111, 25'b1111111111101000110011001, 25'b1111111111001111011001000, 25'b0000000001111100101100011, 25'b1111111111110011011010001, 25'b1111111111010100101001000},
{25'b1111111101100111010110111, 25'b0000000000000110000110001, 25'b1111111101011110111011110, 25'b0000000001101111011010011, 25'b0000000100000111001010001, 25'b0000000000011101101110010, 25'b0000000000000000111110110, 25'b0000000000001100000101001, 25'b1111111111111111111111100, 25'b0000000000100000110000111, 25'b0000000101001101000100101, 25'b1111111111111111111011100, 25'b0000000001100001100101111, 25'b0000000010011111011110010, 25'b0000000011000100110000101, 25'b0000000100001100110101000, 25'b0000000000000000000000110, 25'b1111111110000101100110100, 25'b0000000001010110000101101, 25'b1111111111111110100110000, 25'b1111111101011100101101100, 25'b1111111111000101111011010, 25'b0000000000000011011100110, 25'b1111111111101010110011100, 25'b1111111101111111101010000, 25'b0000000111100000001001000, 25'b1111111111000111110010000, 25'b0000000000000000000000111, 25'b0000000000000000000000110, 25'b0000000011100010000011110, 25'b0000000000010110101100110, 25'b0000000001100100010011000},
{25'b0000000001101100000110100, 25'b1111111111111011000001110, 25'b0000000000000000000100101, 25'b1111111111110100111010001, 25'b0000000000010100111000111, 25'b1111111111110110010000010, 25'b1111111111111111111011101, 25'b0000000000101000001010110, 25'b0000000000110110000111000, 25'b1111111110111001110111001, 25'b0000000000100011110110101, 25'b0000000000101111111110010, 25'b0000000000000011000010010, 25'b0000000001010101001100010, 25'b1111111111000110011000110, 25'b1111111100110011111111000, 25'b0000000000000000000000110, 25'b1111111111111100011011011, 25'b1111111111111001001010111, 25'b1111111110000000010111100, 25'b1111111111111111101101111, 25'b0000000000000000000001100, 25'b1111111111001100000110011, 25'b1111111111111100011000100, 25'b1111111111100111101011111, 25'b0000000000100111111000001, 25'b0000000001011111101010110, 25'b1111111111100001011010100, 25'b1111111111110011011011100, 25'b1111111111110101101100110, 25'b0000000000000110111010111, 25'b1111111110011011100010111},
{25'b1111111111010010100001010, 25'b0000000001100010011010010, 25'b0000000000000000000001111, 25'b0000000000000000000000110, 25'b0000000011001010110101000, 25'b0000000001010010011111100, 25'b1111111111111111111111101, 25'b1111111101110001111001111, 25'b0000000000011110001011010, 25'b1111111101001101011010111, 25'b1111111010011000110011110, 25'b1111111111111111111110111, 25'b0000000000000000000101010, 25'b0000000001101101110100001, 25'b0000000000011100011010010, 25'b0000000000000000000001100, 25'b1111111110101011111010100, 25'b0000000000000000000101111, 25'b0000000000000001101110010, 25'b0000000000001111100001001, 25'b0000000000111110011010100, 25'b1111111111111001011111001, 25'b1111111110100011110011000, 25'b0000000000000010000110111, 25'b1111111111111101000110110, 25'b0000000100010100110110001, 25'b0000000001010011100111011, 25'b1111111111111111111001111, 25'b1111111111101101110111010, 25'b0000000010101011000101101, 25'b1111111111110101110011101, 25'b1111111111101001100101110},
{25'b1111111101111010000111110, 25'b0000000000101100110111111, 25'b1111111111110111000111111, 25'b1111111111111111111110110, 25'b1111111111000000111110100, 25'b1111111110011111010100100, 25'b0000000000001100010011011, 25'b0000000000100100111010111, 25'b1111111111111111111111110, 25'b1111111111010100001011101, 25'b1111111101101101011010110, 25'b0000000000110011011010010, 25'b0000000001001101110111010, 25'b0000000000000000000000100, 25'b0000000011010110110001101, 25'b1111111101110000001100100, 25'b0000000000011010100111010, 25'b1111111110011011111001100, 25'b0000000001001000001100001, 25'b1111111111111111111100100, 25'b1111111111110110001001000, 25'b0000000000010001111111011, 25'b0000000000011111011010000, 25'b0000000000000000000010000, 25'b1111111110000001100111010, 25'b0000000000000111111110000, 25'b1111111101110000111100110, 25'b1111111111110101110100110, 25'b1111111111111111111100100, 25'b0000000010101100111111101, 25'b1111111111001111010101111, 25'b0000000000000000000100100},
{25'b1111111111111111111111000, 25'b0000000000011101011001101, 25'b0000000000000000000100100, 25'b0000000001100100001010111, 25'b1111111111100010000001101, 25'b1111111111110100111110001, 25'b0000000000001110111111010, 25'b1111111111111110100000101, 25'b1111111111110100001001110, 25'b0000000010100100000000100, 25'b0000000010110010111110001, 25'b0000000000000000001011001, 25'b1111111110101010110111110, 25'b1111111101001100001110001, 25'b1111111111110011000001011, 25'b0000000000000000000010100, 25'b0000000000000000000010100, 25'b1111111111101111101100010, 25'b1111111110000110000001011, 25'b0000000001100001111000100, 25'b0000000000000000100010100, 25'b0000000001011110111110010, 25'b1111111111111111111100000, 25'b0000000010001111111111100, 25'b0000000000011111101011100, 25'b0000000001001110011011000, 25'b0000000001110100100111110, 25'b1111111111110010110000101, 25'b1111111110011011110010111, 25'b1111111110001111001100100, 25'b1111111111111110101101001, 25'b1111111101010100110000110},
{25'b1111111111000110000100000, 25'b1111111111111111111111000, 25'b0000000000011110100010011, 25'b1111111110010100110000001, 25'b0000000000010110000011001, 25'b1111111111111111111110010, 25'b1111111111001000011001111, 25'b1111111111111101100010100, 25'b1111111111011111111001100, 25'b0000000000001001100000111, 25'b0000000000010011111101100, 25'b1111111111101101101101111, 25'b0000000000000100001110011, 25'b0000000000110000000010011, 25'b1111111101011111111111011, 25'b1111111111000001010111100, 25'b0000000000111010011010010, 25'b1111111111010010101101111, 25'b0000000000000000000001010, 25'b1111111111111001100100101, 25'b0000000000110001011010000, 25'b0000000000000010000011010, 25'b1111111111111000000010011, 25'b0000000000001010111000010, 25'b0000000001000100111111000, 25'b1111111111100101011001101, 25'b0000000000000000000011000, 25'b1111111110001100010111010, 25'b1111111111001101111001001, 25'b1111111111111110001101010, 25'b0000000000101100011000110, 25'b0000000000000000000101111},
{25'b1111111101111010111100001, 25'b0000000001101011100111100, 25'b1111111111111111111111001, 25'b1111111111111110010011000, 25'b1111111111111101100010000, 25'b0000000000101100111000101, 25'b1111111111111111111100001, 25'b0000000011000101101001110, 25'b1111111111111100001110000, 25'b1111111111111111111111011, 25'b0000000000110100101100001, 25'b0000000000001010011111101, 25'b0000000000000001101010101, 25'b0000000000000000000011110, 25'b0000000000011111001011001, 25'b0000000001010100100001110, 25'b0000000000101101100111000, 25'b0000000000101010101011101, 25'b1111111111111101110100100, 25'b0000000001001110101010000, 25'b0000000000011001110001000, 25'b0000000000001010010111111, 25'b1111111111111101110011000, 25'b0000000001000001000001010, 25'b1111111111100110100000010, 25'b1111111110101001001111101, 25'b1111111111101000010110111, 25'b1111111111111111111111001, 25'b0000000000011010000000110, 25'b0000000000000111100110101, 25'b0000000000110010000001000, 25'b0000000001111010101010010},
{25'b1111111111111011001110000, 25'b1111111110011100010101111, 25'b0000000000001101001110001, 25'b1111111111111111110000001, 25'b0000000011101010100001011, 25'b1111111111001010111010110, 25'b1111111101101101101011011, 25'b0000000000000000000011010, 25'b0000000000000000000010000, 25'b1111111111111001011001011, 25'b0000000000001100011001111, 25'b0000000001101111110011110, 25'b0000000001010010011010111, 25'b0000000000000010101110111, 25'b0000000000001000100010011, 25'b1111111111010011010001010, 25'b0000000000001000100010011, 25'b1111111111110110010010001, 25'b0000000000000000000001101, 25'b0000000000010011010011000, 25'b1111111111110110011010101, 25'b0000000000000100111010000, 25'b0000000001000100001010011, 25'b0000000000001001011100100, 25'b1111111111111100111010100, 25'b1111111110010110010110000, 25'b0000000000110100000001011, 25'b1111111111111111111111000, 25'b1111111111111111111010011, 25'b1111111111100100110010010, 25'b1111111111111010100000100, 25'b1111111111101111111110111},
{25'b0000000000000001110100011, 25'b1111111111101111110011001, 25'b1111111111011111101110010, 25'b1111111111001000000000010, 25'b1111111101110100000100110, 25'b0000000010011100000001001, 25'b0000000000000000000011111, 25'b0000000000101011001111110, 25'b0000000001001001011110000, 25'b0000000000000011010010001, 25'b1111111111110111010101110, 25'b0000000001111001110001100, 25'b0000000000111001010011101, 25'b1111111110100010011010101, 25'b1111111111010110011100000, 25'b1111111111110101011101101, 25'b1111111110011010000000001, 25'b1111111111111011100011101, 25'b0000000000000000000011011, 25'b1111111111111110110101001, 25'b0000000000100111111011101, 25'b1111111111011100111111101, 25'b0000000000000000000000110, 25'b0000000000010011101101001, 25'b1111111111111111111110101, 25'b1111111110101000100001101, 25'b0000000000101000000111101, 25'b0000000000000000000110101, 25'b0000000000001011011100000, 25'b0000000000000010110011101, 25'b1111111110101111000101101, 25'b0000000000000101010100011},
{25'b1111111111001101110011101, 25'b1111111111010111101101110, 25'b0000000000010011100100010, 25'b1111111111100000001110101, 25'b1111111111101001000000011, 25'b0000000000011101101111101, 25'b1111111111111110101100001, 25'b0000000000001000111100011, 25'b0000000000100001100010001, 25'b1111111111111111111010001, 25'b0000000000011111101011100, 25'b1111111111011111011010100, 25'b1111111111111101100001000, 25'b1111111111111111111101000, 25'b0000000000011010011110101, 25'b1111111111111111111110101, 25'b0000000001111101000011100, 25'b1111111111111011100011111, 25'b0000000000111111100000000, 25'b1111111111010100100010110, 25'b0000000000101000100000110, 25'b0000000000010000000101100, 25'b0000000000010101100110101, 25'b0000000000001001010010011, 25'b1111111111101011001010010, 25'b1111111110111000101000011, 25'b1111111110111101101011100, 25'b0000000000011011101000000, 25'b1111111111101010100100110, 25'b0000000000000000001001011, 25'b1111111111111000111111010, 25'b0000000000111011011010101},
{25'b1111111111111111111110100, 25'b1111111110011000010111010, 25'b1111111110011010011111001, 25'b1111111111111111111110011, 25'b0000000010100001101000000, 25'b1111111111101000110001000, 25'b0000000000000000000010101, 25'b0000000001111011101110011, 25'b1111111111011010001111101, 25'b0000000000000000000001001, 25'b1111111110010101000100011, 25'b1111111110000010100001100, 25'b0000000001110010110000110, 25'b0000000000100110101100011, 25'b1111111111100000111100100, 25'b1111111110111001111011011, 25'b0000000000101100001000101, 25'b0000000000000000000111011, 25'b1111111111000011001001001, 25'b0000000000000110110011010, 25'b0000000000010001110011001, 25'b1111111111101001010111101, 25'b0000000001001000101101011, 25'b1111111100000101001100110, 25'b0000000000001010011111110, 25'b0000000000111101001100110, 25'b1111111111110101011101111, 25'b0000000000000011110100010, 25'b1111111111000100010010010, 25'b1111111111111111111101101, 25'b1111111111001100100000001, 25'b1111111111111001110101011},
{25'b0000000000110110011011100, 25'b0000000001011000010111100, 25'b0000000010001100111111111, 25'b1111111111001011101001011, 25'b0000000001101010100001011, 25'b0000000001001110011011000, 25'b0000000000000000001000001, 25'b0000000001110100100110001, 25'b0000000001011011011011111, 25'b1111111111100100101001110, 25'b0000000010110011100111101, 25'b1111111110100110100110101, 25'b0000000010011111000100010, 25'b0000000001110010010001100, 25'b1111111011101101010100011, 25'b1111111111111111110000001, 25'b0000000000000000000001000, 25'b0000000000000001011110011, 25'b0000000001000010100010101, 25'b1111111101111111001011110, 25'b0000000000111000101111111, 25'b1111111111001001110000000, 25'b1111111110000010011111100, 25'b1111111111010111110110001, 25'b0000000001010100010100011, 25'b1111111101010111000110011, 25'b1111111110101011100101010, 25'b1111111111110101011101001, 25'b1111111111111111111101100, 25'b1111111101101111100010110, 25'b0000000001100101001111101, 25'b0000000000000000000110010},
{25'b1111111111110011011000011, 25'b0000000000000000001011110, 25'b1111111111111111111111010, 25'b1111111111111111111111101, 25'b1111111110100110000110101, 25'b0000000000000010010110101, 25'b0000000000000010000111001, 25'b1111111111111100001010000, 25'b1111111111111001110011111, 25'b1111111111110100001111000, 25'b0000000000100011100101001, 25'b1111111111111111110100000, 25'b0000000000010101001110101, 25'b1111111110101000011001110, 25'b0000000000011011010111111, 25'b1111111111111111110100011, 25'b0000000000100100000001101, 25'b0000000001110010100110111, 25'b1111111110100101101101011, 25'b0000000000001101010010010, 25'b1111111111100110101001000, 25'b0000000000100000111011101, 25'b0000000000110000101011000, 25'b1111111111101010001011001, 25'b1111111110111111101100010, 25'b0000000000000101010001011, 25'b0000000011010100010011011, 25'b1111111111111001110011100, 25'b1111111111111100000101101, 25'b0000000001010011000001101, 25'b0000000000000000000011011, 25'b0000000011011100101011100},
{25'b1111111101111010011110011, 25'b0000000000001001010000011, 25'b1111111111001000100111110, 25'b0000000001100010000010000, 25'b0000000000011100000101101, 25'b1111111111110111111010001, 25'b1111111111111111111111100, 25'b1111111111111111111111111, 25'b1111111110110010011001111, 25'b1111111111110111100011110, 25'b0000000000000000000010011, 25'b1111111101110001110110011, 25'b0000000000000011001101011, 25'b1111111111110101110100101, 25'b1111111111111111011000000, 25'b1111111111111111111101000, 25'b1111111111100010001000101, 25'b0000000000000001011001001, 25'b0000000000000000110011110, 25'b0000000000101000101000000, 25'b0000000000000100011111001, 25'b0000000000000000000000100, 25'b0000000000000000000010010, 25'b1111111111111101111011100, 25'b0000000000000000000100110, 25'b0000000000000100101100000, 25'b0000000010010100110101000, 25'b1111111111111111111111100, 25'b1111111111111111111101001, 25'b1111111111110101100100101, 25'b0000000000101100110100010, 25'b1111111111111001011110101},
{25'b1111111111111111100110001, 25'b1111111111011001010000001, 25'b0000000000110100010011010, 25'b0000000000001010001110110, 25'b1111111110100000110101110, 25'b0000000000000000001010000, 25'b0000000001001001001101000, 25'b1111111111111111111101101, 25'b0000000000000000000000111, 25'b1111111111100110110000101, 25'b0000000000011101011011111, 25'b0000000000000100110111011, 25'b0000000001010010110101011, 25'b1111111101110011101001110, 25'b1111111111100111110011101, 25'b1111111111111011100110010, 25'b0000000000110111010101110, 25'b1111111110011101101011101, 25'b0000000000000101011100000, 25'b1111111100111110110100010, 25'b1111111111111011001010101, 25'b1111111111100001100011100, 25'b1111111111110101101011100, 25'b0000000001001011101100100, 25'b1111111111101100111011100, 25'b1111111110111000000011101, 25'b0000000000010111001000011, 25'b0000000000000000000101001, 25'b0000000001100101010101010, 25'b0000000010000101111101000, 25'b1111111110101100000001000, 25'b1111111110001101000000001},
{25'b0000000000010001010001001, 25'b0000000000000110100010011, 25'b1111111110010101111111100, 25'b1111111111110001011110000, 25'b1111111111111111111110010, 25'b0000000000000000100011110, 25'b0000000000011011001101000, 25'b0000000001101001010011110, 25'b0000000000000000000001010, 25'b0000000000000101001100100, 25'b0000000000010001111011011, 25'b1111111101110101111010110, 25'b1111111111101110111101001, 25'b1111111101100101011100010, 25'b0000000001111011000110000, 25'b0000000000000000000110101, 25'b1111111111111111110011011, 25'b1111111101011011111101100, 25'b1111111111111111111011110, 25'b1111111111101100111101000, 25'b1111111111111010101011001, 25'b0000000000000000000000010, 25'b0000000000001111111101111, 25'b1111111111011001100001101, 25'b0000000000001101100110111, 25'b0000000001101001001100000, 25'b0000000001101101001010100, 25'b0000000001100011111111001, 25'b0000000001001110110110111, 25'b0000000000000000000011001, 25'b0000000000011101001111100, 25'b0000000011001000100101100},
{25'b1111111111111001100010111, 25'b1111111111000011000111101, 25'b0000000001100011101011011, 25'b1111111111100101101010101, 25'b0000000000010001110111011, 25'b0000000000101010111110011, 25'b1111111111111111111111111, 25'b1111111110110110100010101, 25'b1111111111101010001100011, 25'b1111111101100110001101111, 25'b0000000001110010100000101, 25'b0000000000000000111110010, 25'b0000000001101011010010001, 25'b0000000010101011100011011, 25'b1111111111100010001100111, 25'b1111111100100001000111100, 25'b1111111111100101011010101, 25'b0000000001111000010010111, 25'b1111111110110111100101111, 25'b1111111111001010100101110, 25'b0000000000001111001101101, 25'b0000000000000000010000001, 25'b1111111101110100011110110, 25'b1111111111001111000010100, 25'b1111111111110101111100110, 25'b1111111111100000110100010, 25'b0000000000011100101111101, 25'b0000000010110100001000000, 25'b0000000000111110110110100, 25'b1111111111111111111110100, 25'b0000000000010100101010111, 25'b0000000000000111000100111},
{25'b0000000000001010110111011, 25'b0000000001110100001001110, 25'b0000000000000000000001111, 25'b0000000001001011101001110, 25'b0000000011010100110011101, 25'b1111111111010100010010111, 25'b1111111111111111111111000, 25'b1111111111110100101010110, 25'b0000000001001011000000101, 25'b1111111111001110111110011, 25'b1111111111111111101010111, 25'b0000000001010101010101001, 25'b0000000000000010001011011, 25'b0000000000000111000001100, 25'b1111111001111001000101001, 25'b1111111111101011101011001, 25'b0000000000000000000000001, 25'b0000000000110011011000000, 25'b1111111111111111001001000, 25'b0000000001001100011100101, 25'b1111111111111111111100011, 25'b1111111111010011110001101, 25'b1111111101110000001010000, 25'b0000000000100001011111101, 25'b0000000001001001001100001, 25'b1111111011100100000100000, 25'b1111111111111111111100101, 25'b0000000000000000000010111, 25'b0000000010001011010010111, 25'b1111111100110010110110111, 25'b0000000000000000011101101, 25'b1111111111111110011100011},
{25'b0000000000000010011010100, 25'b1111111110101001000011111, 25'b0000000000001101110100010, 25'b1111111111111100001011011, 25'b0000000000001101010101001, 25'b0000000010000111011100011, 25'b1111111101000110011101110, 25'b0000000000001000110011110, 25'b0000000001101100011001011, 25'b1111111110101001101011010, 25'b1111111111111010000011110, 25'b0000000000001100100001001, 25'b1111111111111101101101110, 25'b0000000000101101110010110, 25'b0000000000011011011111001, 25'b1111111111111011101111101, 25'b0000000000010001001010111, 25'b0000000000000000000100111, 25'b0000000000000101100010000, 25'b0000000001100001001111111, 25'b1111111111111000110100010, 25'b1111111110000100000000001, 25'b1111111101100101001001111, 25'b1111111111001110011010100, 25'b1111111101101000110010011, 25'b0000000000110101010000010, 25'b0000000010011111100011010, 25'b0000000001011110011000011, 25'b1111111111111101010101010, 25'b1111111110100000100111001, 25'b1111111110110000011100111, 25'b0000000000001111010010111},
{25'b0000000000001101010010110, 25'b1111111110000101101110110, 25'b1111111111111011101011010, 25'b0000000000100110100001101, 25'b1111111110000101100000110, 25'b0000000000101011011100111, 25'b1111111111111111111110000, 25'b1111111111111111111101011, 25'b1111111111111111111111011, 25'b0000000000000000000011101, 25'b0000000001000011101011101, 25'b1111111111111011100101100, 25'b0000000000000010011111110, 25'b0000000000000000000100001, 25'b0000000000100000100110110, 25'b1111111111111011101011111, 25'b0000000000000000101101001, 25'b1111111111111111110101000, 25'b1111111110101101100011111, 25'b1111111101111110100011100, 25'b1111111111111111110110100, 25'b1111111101110111010101001, 25'b1111111110110010111001110, 25'b1111111110100000110101011, 25'b0000000011100011111111011, 25'b0000000000000100100000001, 25'b1111111111110100001101111, 25'b0000000001010001001111011, 25'b0000000011100101110000000, 25'b0000000001100101000101101, 25'b1111111011110000100001100, 25'b1111111111010000100000111},
{25'b0000000001100000001110011, 25'b1111111111111111111001110, 25'b0000000001000000010000111, 25'b1111111111111010111010101, 25'b0000000001111011110101111, 25'b1111111111011011011111110, 25'b0000000000010010001000011, 25'b0000000001101011000100010, 25'b0000000001000100100011100, 25'b1111111101111010010100011, 25'b1111111111110000010000000, 25'b0000000000011111011101000, 25'b0000000000010001101001110, 25'b1111111111111100010000110, 25'b0000000000010101101111001, 25'b0000000000000000000100010, 25'b0000000001011100110001001, 25'b0000000000001000111110100, 25'b0000000001011111110010111, 25'b1111111111101111001110111, 25'b1111111111011111011001111, 25'b1111111111101100110110011, 25'b1111111111111111111100010, 25'b0000000001001101010001110, 25'b1111111111001100001100110, 25'b1111111111111110011010011, 25'b0000000000000000000000001, 25'b0000000000000000000100010, 25'b0000000000000000000010000, 25'b0000000001001010110001110, 25'b1111111110101101111010001, 25'b1111111111111010000011101},
{25'b1111111111111111110101100, 25'b1111111111111000000110010, 25'b1111111110001000111100011, 25'b0000000001001000110101011, 25'b0000000000111001001000010, 25'b1111111111100011111100111, 25'b1111111111111111111101111, 25'b1111111111000101111010001, 25'b0000000000000001101110010, 25'b1111111111111111111010101, 25'b1111111110110010110110011, 25'b1111111111000000111100010, 25'b0000000001111010101000100, 25'b0000000000000000000000001, 25'b1111111111011111010011000, 25'b1111111111111111111111001, 25'b0000000000110110110011100, 25'b1111111111111111111101011, 25'b1111111111111111111111110, 25'b1111111111001000101101101, 25'b0000000001010000111110101, 25'b0000000000000000000001001, 25'b0000000000100111111111000, 25'b1111111111111000101011000, 25'b0000000000101000001100010, 25'b0000000000000000100100001, 25'b0000000000000000000001110, 25'b0000000000111101101000100, 25'b1111111111001110110100110, 25'b1111111111110100001101010, 25'b0000000000101001000110110, 25'b1111111111100100111001101},
{25'b1111111111111011101110000, 25'b1111111110110001000000100, 25'b0000000010011000001010110, 25'b1111111111101111010111111, 25'b0000000000110010010001111, 25'b1111111110110110110001000, 25'b0000000000000000000001001, 25'b0000000000001000110000000, 25'b1111111110000101010111101, 25'b1111111111111100101110100, 25'b1111111111100000010100011, 25'b0000000000001110111001001, 25'b1111111110101100000011111, 25'b0000000000100011010011010, 25'b0000000000110011110010001, 25'b0000000000011100000011011, 25'b0000000000010101111101110, 25'b1111111111110110010000110, 25'b1111111101001010101101011, 25'b1111111111111100100011010, 25'b1111111111110001011011101, 25'b0000000000100011110011010, 25'b1111111111100011100100010, 25'b1111111111111111111111111, 25'b0000000000110010100111011, 25'b1111111111110100010101110, 25'b1111111111111100010011010, 25'b0000000001100011100101101, 25'b1111111110011010000111000, 25'b1111111110110100011100001, 25'b0000000001011001110011111, 25'b0000000000001001001100011},
{25'b0000000001101110010100101, 25'b0000000000110011100010001, 25'b0000000000000000001100100, 25'b1111111111010111010011100, 25'b1111111111101011111010010, 25'b1111111111111111110010010, 25'b0000000000000000000001001, 25'b1111111111101110010011011, 25'b1111111111100000001101010, 25'b1111111111100001101010101, 25'b0000000000000000000101011, 25'b0000000000101000100010111, 25'b0000000000000001101000110, 25'b0000000000001101100010000, 25'b1111111111110100100100100, 25'b0000000000000001011110100, 25'b1111111111011000101111010, 25'b0000000000000000001001110, 25'b1111111111111011100000000, 25'b1111111111111111110110011, 25'b0000000000000000100110011, 25'b0000000000001111001101110, 25'b0000000000011000111000011, 25'b0000000000000000000001100, 25'b0000000000000000000100100, 25'b1111111101100011101101111, 25'b1111111111001100111111010, 25'b0000000000000001101100010, 25'b0000000000000101001111010, 25'b0000000000000000010101110, 25'b1111111111010010101010011, 25'b0000000000000101100000000},
{25'b0000000000110000000010010, 25'b1111111011110100100110011, 25'b1111111111111111111110100, 25'b1111111111101100101111101, 25'b1111111111000100011000101, 25'b1111111111111101100010111, 25'b0000000000000000000000110, 25'b0000000010001100001111010, 25'b1111111111110100110010000, 25'b1111111111111010011000001, 25'b0000000000010101001000000, 25'b1111111101010110110111010, 25'b0000000000000110001001001, 25'b1111111110001111110000010, 25'b0000000010111000111100100, 25'b1111111111110010100111101, 25'b1111111111000110000001100, 25'b1111111101110011111101110, 25'b1111111111111101010011101, 25'b1111111101001010110011011, 25'b1111111100110000101110000, 25'b1111111111111111111011100, 25'b0000000000000000000111011, 25'b0000000000000000000001001, 25'b0000000000111110011110010, 25'b1111111111111100011011111, 25'b1111111110110011101010011, 25'b1111111111101101011001010, 25'b1111111111111010000010001, 25'b0000000000000000000011110, 25'b1111111111110111111000110, 25'b1111111101001100110100001}
};
localparam logic signed [24:0] bias [32] = '{
25'b0000000001000011100110001,
25'b0000000001101011101101000,
25'b0000000000110010111011000,
25'b0000000000110100100011101,
25'b1111111000101011110011111,
25'b1111111110001101000101010,
25'b0000000011011010010001000,
25'b1111111101011100100110110,
25'b1111111110110101010001101,
25'b0000000101011001100011110,
25'b0000000000011011110010010,
25'b0000000001110000110100111,
25'b1111111010101110110011110,
25'b1111111100001111101101001,
25'b0000000011010100110011110,
25'b0000000101011111011111000,
25'b1111111111000010110001001,
25'b0000000011011001011010001,
25'b0000000001101101011011010,
25'b0000000010000000100101100,
25'b0000000010110101101110110,
25'b0000000001101010100011100,
25'b0000000001000101100011101,
25'b0000000001110110110000000,
25'b1111111111010100001001011,
25'b1111111110111000011111000,
25'b1111111110110000100001111,
25'b1111111101011100001000001,
25'b0000000000000111100110101,
25'b1111111110010110110111101,
25'b0000000001110000011011111,
25'b1111111110000110011100000
};
endpackage