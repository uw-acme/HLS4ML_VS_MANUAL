// Width: 27
// NFRAC: 13
package dense_3_27_14;

localparam logic signed [26:0] weights [32][32] = '{ 
{27'b111111111111111111001101101, 27'b111111111111111001000000010, 27'b111111111111111001100000100, 27'b111111111111111100111100111, 27'b000000000000000101011111011, 27'b000000000000000000101100111, 27'b111111111111111111110010111, 27'b111111111111111111111111001, 27'b111111111111111111111111111, 27'b111111111111111111111111110, 27'b000000000000000010000001000, 27'b111111111111110111100100011, 27'b111111111111111111000010111, 27'b000000000000001101100011011, 27'b111111111111111100001000101, 27'b111111111111110001000100111, 27'b111111111111111111011010110, 27'b000000000000000001110010000, 27'b000000000000000110111101011, 27'b111111111111111010011011010, 27'b111111111111101110111100110, 27'b111111111111111111010000111, 27'b000000000000000000110010011, 27'b111111111111111001100011000, 27'b000000000000000000000000001, 27'b000000000000010000001100111, 27'b111111111111101000101100100, 27'b111111111111111100011101000, 27'b111111111111111001110010001, 27'b111111111111111101100110010, 27'b000000000000000110110001001, 27'b111111111111111101011100110}, 
{27'b000000000000001011111101101, 27'b000000000000011011101011100, 27'b000000000000000110011011101, 27'b111111111111110101011110100, 27'b000000000000000011111010001, 27'b111111111111111011101000000, 27'b111111111111111110010000111, 27'b000000000000010001011100000, 27'b000000000000000000000110000, 27'b111111111111111111111111111, 27'b111111111111111111011111011, 27'b111111111111110110100101101, 27'b111111111111111100110001110, 27'b000000000000001000101001010, 27'b111111111111011110010011101, 27'b111111111111111000011101011, 27'b111111111111111111111111111, 27'b111111111111111111110111100, 27'b111111111111111111001010000, 27'b111111111111111101010111110, 27'b111111111111111011110111011, 27'b111111111111111011100110000, 27'b000000000000000000010001101, 27'b111111111111111111111110010, 27'b111111111111111111111001011, 27'b111111111111101110110110001, 27'b000000000000000000001100000, 27'b000000000000000111100010010, 27'b111111111111111110111111001, 27'b111111111111110100111101101, 27'b000000000000000000000010110, 27'b000000000000000000100110110}, 
{27'b111111111111110000001111001, 27'b000000000000000010111100100, 27'b000000000000000000001010111, 27'b000000000000000101001010011, 27'b111111111111110101111010100, 27'b000000000000000000000000100, 27'b000000000000000000000001101, 27'b111111111111110010100100101, 27'b000000000000001000100100110, 27'b111111111111111011110011101, 27'b111111111111111011110110010, 27'b111111111111101000001101011, 27'b111111111111111011000001100, 27'b000000000000001000001011001, 27'b000000000000000100001110001, 27'b111111111111111111111110010, 27'b111111111111111110001010111, 27'b111111111111111111100111110, 27'b111111111111110010111101111, 27'b000000000000000000000011001, 27'b000000000000000001111111101, 27'b000000000000000001000110101, 27'b000000000000000011010110001, 27'b000000000000001110000101001, 27'b000000000000000000100110110, 27'b111111111111110011011000111, 27'b000000000000001100010001110, 27'b000000000000000000000000101, 27'b000000000000000010101001110, 27'b111111111111111111101001011, 27'b000000000000000000000000111, 27'b000000000000100100010011010}, 
{27'b000000000000001101011001110, 27'b111111111111111111111111111, 27'b111111111111111100111000111, 27'b000000000000010100111100000, 27'b000000000000010011101001100, 27'b000000000000000000000000010, 27'b000000000000000001001011011, 27'b000000000000001101000001010, 27'b111111111111111001101010100, 27'b111111111111111111111111110, 27'b111111111111110010110100111, 27'b000000000000000001111010100, 27'b000000000000000100010000111, 27'b111111111111110100000010101, 27'b000000000000000001011111110, 27'b111111111111111101011100010, 27'b111111111111111111111111110, 27'b111111111111111010001011001, 27'b000000000000000000100111011, 27'b000000000000000000111000100, 27'b000000000000000000010000010, 27'b111111111111111110110101010, 27'b000000000000010011000110010, 27'b000000000000001010111110001, 27'b000000000000001010100010100, 27'b000000000000000111111100010, 27'b000000000000001010111011100, 27'b000000000000000000000000011, 27'b111111111111111110000111001, 27'b000000000000001110011111111, 27'b000000000000000111111111000, 27'b111111111111111101001100001}, 
{27'b000000000000010000000000100, 27'b111111111111111110100000010, 27'b111111111111110100111010001, 27'b111111111111100111111100110, 27'b000000000000001111010001110, 27'b000000000000000000000000010, 27'b111111111111110010110111111, 27'b111111111111110110111101001, 27'b111111111111111110100000101, 27'b111111111111100110000110101, 27'b111111111111011100101001010, 27'b000000000000001111001000000, 27'b000000000000010101011001101, 27'b000000000000010000101111110, 27'b111111111111101101100110010, 27'b111111111111100111001100110, 27'b000000000000000000000000001, 27'b111111111111111011011110011, 27'b000000000000000110011011000, 27'b000000000000000100011100000, 27'b111111111111111001111110001, 27'b111111111111111111110010111, 27'b000000000000010111000101111, 27'b111111111111010100000000100, 27'b000000000000000010110100010, 27'b111111111111101010111011010, 27'b000000000000000010000110001, 27'b111111111111111000000011110, 27'b111111111111110110011100110, 27'b111111111111111111111111010, 27'b000000000000000010001111010, 27'b000000000000010010100100111}, 
{27'b000000000000000001011000011, 27'b111111111111111110101011010, 27'b111111111111110110001011001, 27'b111111111111110111101010111, 27'b000000000000001011111001010, 27'b000000000000000000000000010, 27'b111111111111110111000011000, 27'b111111111111111011101001001, 27'b111111111111110010010011001, 27'b111111111111111101111100110, 27'b111111111111111111111111000, 27'b000000000000000101001000010, 27'b000000000000000000000000000, 27'b000000000000001011011100101, 27'b111111111111101111110100001, 27'b111111111111111011111010100, 27'b000000000000000010110110011, 27'b111111111111110110100111111, 27'b111111111111111001101011011, 27'b111111111111111111111111110, 27'b000000000000000000011000111, 27'b000000000000001001100101101, 27'b000000000000001110111100011, 27'b111111111111111111101010001, 27'b111111111111111111111111001, 27'b000000000000001100110100101, 27'b111111111111101110011010100, 27'b111111111111111111111111110, 27'b111111111111111000011011100, 27'b111111111111111110110100100, 27'b111111111111111111111001100, 27'b000000000000000000001101010}, 
{27'b000000000000000010000101010, 27'b111111111111110101010111001, 27'b000000000000000011011101111, 27'b111111111111111110110001001, 27'b111111111111111111110000100, 27'b000000000000000100110110000, 27'b111111111111111100100110111, 27'b111111111111101010010101010, 27'b111111111111111111111111110, 27'b111111111111111001010101010, 27'b111111111111110001011000100, 27'b000000000000001111000111000, 27'b000000000000000000001110100, 27'b000000000000010101111001100, 27'b000000000000011010100001001, 27'b000000000000000000000101010, 27'b111111111111111111111111111, 27'b111111111111110101111010010, 27'b111111111111111110000001001, 27'b000000000000001000101111110, 27'b111111111111100111111111110, 27'b000000000000000100111111011, 27'b000000000000001010011100010, 27'b000000000000000000100110111, 27'b000000000000000100110011011, 27'b000000000000100111110010010, 27'b111111111111110011011000110, 27'b111111111111111101000110011, 27'b111111111111111001111011001, 27'b000000000000001111100101100, 27'b111111111111111110011011010, 27'b111111111111111010100101001}, 
{27'b111111111111101100111010110, 27'b000000000000000000110000110, 27'b111111111111101011110111011, 27'b000000000000001101111011010, 27'b000000000000100000111001010, 27'b000000000000000011101101110, 27'b000000000000000000000111110, 27'b000000000000000001100000101, 27'b111111111111111111111111111, 27'b000000000000000100000110000, 27'b000000000000101001101000100, 27'b111111111111111111111111011, 27'b000000000000001100001100101, 27'b000000000000010011111011110, 27'b000000000000011000100110000, 27'b000000000000100001100110101, 27'b000000000000000000000000000, 27'b111111111111110000101100110, 27'b000000000000001010110000101, 27'b111111111111111111110100110, 27'b111111111111101011100101101, 27'b111111111111111000101111011, 27'b000000000000000000011011100, 27'b111111111111111101010110011, 27'b111111111111101111111101010, 27'b000000000000111100000001000, 27'b111111111111111000111110010, 27'b000000000000000000000000000, 27'b000000000000000000000000000, 27'b000000000000011100010000011, 27'b000000000000000010110101100, 27'b000000000000001100100010010}, 
{27'b000000000000001101100000110, 27'b111111111111111111011000001, 27'b000000000000000000000000100, 27'b111111111111111110100111010, 27'b000000000000000010100111000, 27'b111111111111111110110010000, 27'b111111111111111111111111011, 27'b000000000000000101000001010, 27'b000000000000000110110000111, 27'b111111111111110111001110111, 27'b000000000000000100011110110, 27'b000000000000000101111111110, 27'b000000000000000000011000010, 27'b000000000000001010101001100, 27'b111111111111111000110011000, 27'b111111111111100110011111110, 27'b000000000000000000000000000, 27'b111111111111111111100011011, 27'b111111111111111111001001010, 27'b111111111111110000000010111, 27'b111111111111111111111101101, 27'b000000000000000000000000001, 27'b111111111111111001100000110, 27'b111111111111111111100011000, 27'b111111111111111100111101011, 27'b000000000000000100111111000, 27'b000000000000001011111101010, 27'b111111111111111100001011010, 27'b111111111111111110011011011, 27'b111111111111111110101101100, 27'b000000000000000000110111010, 27'b111111111111110011011100010}, 
{27'b111111111111111010010100001, 27'b000000000000001100010011010, 27'b000000000000000000000000001, 27'b000000000000000000000000000, 27'b000000000000011001010110101, 27'b000000000000001010010011111, 27'b111111111111111111111111111, 27'b111111111111101110001111001, 27'b000000000000000011110001011, 27'b111111111111101001101011010, 27'b111111111111010011000110011, 27'b111111111111111111111111110, 27'b000000000000000000000000101, 27'b000000000000001101101110100, 27'b000000000000000011100011010, 27'b000000000000000000000000001, 27'b111111111111110101011111010, 27'b000000000000000000000000101, 27'b000000000000000000001101110, 27'b000000000000000001111100001, 27'b000000000000000111110011010, 27'b111111111111111111001011111, 27'b111111111111110100011110010, 27'b000000000000000000010000110, 27'b111111111111111111101000110, 27'b000000000000100010100110110, 27'b000000000000001010011100111, 27'b111111111111111111111111001, 27'b111111111111111101101110111, 27'b000000000000010101011000101, 27'b111111111111111110101110011, 27'b111111111111111101001100101}, 
{27'b111111111111101111010000111, 27'b000000000000000101100110111, 27'b111111111111111110111000111, 27'b111111111111111111111111110, 27'b111111111111111000000111110, 27'b111111111111110011111010100, 27'b000000000000000001100010011, 27'b000000000000000100100111010, 27'b111111111111111111111111111, 27'b111111111111111010100001011, 27'b111111111111101101101011010, 27'b000000000000000110011011010, 27'b000000000000001001101110111, 27'b000000000000000000000000000, 27'b000000000000011010110110001, 27'b111111111111101110000001100, 27'b000000000000000011010100111, 27'b111111111111110011011111001, 27'b000000000000001001000001100, 27'b111111111111111111111111100, 27'b111111111111111110110001000, 27'b000000000000000010001111111, 27'b000000000000000011111011010, 27'b000000000000000000000000010, 27'b111111111111110000001100111, 27'b000000000000000000111111101, 27'b111111111111101110000111100, 27'b111111111111111110101110100, 27'b111111111111111111111111100, 27'b000000000000010101100111111, 27'b111111111111111001111010101, 27'b000000000000000000000000100}, 
{27'b111111111111111111111111110, 27'b000000000000000011101011001, 27'b000000000000000000000000100, 27'b000000000000001100100001010, 27'b111111111111111100010000001, 27'b111111111111111110100111110, 27'b000000000000000001110111111, 27'b111111111111111111110100000, 27'b111111111111111110100001001, 27'b000000000000010100100000000, 27'b000000000000010110010111110, 27'b000000000000000000000001011, 27'b111111111111110101010110111, 27'b111111111111101001100001110, 27'b111111111111111110011000001, 27'b000000000000000000000000010, 27'b000000000000000000000000010, 27'b111111111111111101111101100, 27'b111111111111110000110000001, 27'b000000000000001100001111000, 27'b000000000000000000000100010, 27'b000000000000001011110111110, 27'b111111111111111111111111100, 27'b000000000000010001111111111, 27'b000000000000000011111101011, 27'b000000000000001001110011011, 27'b000000000000001110100100111, 27'b111111111111111110010110000, 27'b111111111111110011011110010, 27'b111111111111110001111001100, 27'b111111111111111111110101101, 27'b111111111111101010100110000}, 
{27'b111111111111111000110000011, 27'b111111111111111111111111111, 27'b000000000000000011110100010, 27'b111111111111110010100110000, 27'b000000000000000010110000011, 27'b111111111111111111111111110, 27'b111111111111111001000011001, 27'b111111111111111111101100010, 27'b111111111111111011111111001, 27'b000000000000000001001100000, 27'b000000000000000010011111101, 27'b111111111111111101101101101, 27'b000000000000000000100001110, 27'b000000000000000110000000010, 27'b111111111111101011111111111, 27'b111111111111111000001010111, 27'b000000000000000111010011010, 27'b111111111111111010010101101, 27'b000000000000000000000000001, 27'b111111111111111111001100100, 27'b000000000000000110001011001, 27'b000000000000000000010000011, 27'b111111111111111111000000010, 27'b000000000000000001010111000, 27'b000000000000001000100111110, 27'b111111111111111100101011001, 27'b000000000000000000000000011, 27'b111111111111110001100010111, 27'b111111111111111001101111001, 27'b111111111111111111110001101, 27'b000000000000000101100011000, 27'b000000000000000000000000101}, 
{27'b111111111111101111010111100, 27'b000000000000001101011100111, 27'b111111111111111111111111111, 27'b111111111111111111110010010, 27'b111111111111111111101100010, 27'b000000000000000101100111000, 27'b111111111111111111111111100, 27'b000000000000011000101101001, 27'b111111111111111111100001101, 27'b111111111111111111111111111, 27'b000000000000000110100101100, 27'b000000000000000001010011111, 27'b000000000000000000001101010, 27'b000000000000000000000000011, 27'b000000000000000011111001011, 27'b000000000000001010100100001, 27'b000000000000000101101100111, 27'b000000000000000101010101011, 27'b111111111111111111101110100, 27'b000000000000001001110101001, 27'b000000000000000011001110001, 27'b000000000000000001010010111, 27'b111111111111111111101110011, 27'b000000000000001000001000001, 27'b111111111111111100110100000, 27'b111111111111110101001001111, 27'b111111111111111101000010110, 27'b111111111111111111111111111, 27'b000000000000000011010000000, 27'b000000000000000000111100110, 27'b000000000000000110010000001, 27'b000000000000001111010101010}, 
{27'b111111111111111111011001110, 27'b111111111111110011100010101, 27'b000000000000000001101001110, 27'b111111111111111111111110000, 27'b000000000000011101010100001, 27'b111111111111111001010111010, 27'b111111111111101101101101011, 27'b000000000000000000000000011, 27'b000000000000000000000000001, 27'b111111111111111111001011001, 27'b000000000000000001100011001, 27'b000000000000001101111110011, 27'b000000000000001010010011010, 27'b000000000000000000010101110, 27'b000000000000000001000100010, 27'b111111111111111010011010001, 27'b000000000000000001000100010, 27'b111111111111111110110010010, 27'b000000000000000000000000001, 27'b000000000000000010011010011, 27'b111111111111111110110011010, 27'b000000000000000000100111001, 27'b000000000000001000100001010, 27'b000000000000000001001011100, 27'b111111111111111111100111010, 27'b111111111111110010110010110, 27'b000000000000000110100000001, 27'b111111111111111111111111110, 27'b111111111111111111111111010, 27'b111111111111111100100110010, 27'b111111111111111111010100000, 27'b111111111111111101111111110}, 
{27'b000000000000000000001110100, 27'b111111111111111101111110011, 27'b111111111111111011111101110, 27'b111111111111111001000000000, 27'b111111111111101110100000100, 27'b000000000000010011100000001, 27'b000000000000000000000000011, 27'b000000000000000101011001111, 27'b000000000000001001001011110, 27'b000000000000000000011010010, 27'b111111111111111110111010101, 27'b000000000000001111001110001, 27'b000000000000000111001010011, 27'b111111111111110100010011010, 27'b111111111111111010110011100, 27'b111111111111111110101011101, 27'b111111111111110011010000000, 27'b111111111111111111011100011, 27'b000000000000000000000000011, 27'b111111111111111111110110101, 27'b000000000000000100111111011, 27'b111111111111111011100111111, 27'b000000000000000000000000000, 27'b000000000000000010011101101, 27'b111111111111111111111111110, 27'b111111111111110101000100001, 27'b000000000000000101000000111, 27'b000000000000000000000000110, 27'b000000000000000001011011011, 27'b000000000000000000010110011, 27'b111111111111110101111000101, 27'b000000000000000000101010100}, 
{27'b111111111111111001101110011, 27'b111111111111111010111101101, 27'b000000000000000010011100100, 27'b111111111111111100000001110, 27'b111111111111111101001000000, 27'b000000000000000011101101111, 27'b111111111111111111110101100, 27'b000000000000000001000111100, 27'b000000000000000100001100010, 27'b111111111111111111111111010, 27'b000000000000000011111101011, 27'b111111111111111011111011010, 27'b111111111111111111101100001, 27'b111111111111111111111111101, 27'b000000000000000011010011110, 27'b111111111111111111111111110, 27'b000000000000001111101000011, 27'b111111111111111111011100011, 27'b000000000000000111111100000, 27'b111111111111111010100100010, 27'b000000000000000101000100000, 27'b000000000000000010000000101, 27'b000000000000000010101100110, 27'b000000000000000001001010010, 27'b111111111111111101011001010, 27'b111111111111110111000101000, 27'b111111111111110111101101011, 27'b000000000000000011011101000, 27'b111111111111111101010100100, 27'b000000000000000000000001001, 27'b111111111111111111000111111, 27'b000000000000000111011011010}, 
{27'b111111111111111111111111110, 27'b111111111111110011000010111, 27'b111111111111110011010011111, 27'b111111111111111111111111110, 27'b000000000000010100001100111, 27'b111111111111111101000110001, 27'b000000000000000000000000010, 27'b000000000000001111011101110, 27'b111111111111111011010001111, 27'b000000000000000000000000001, 27'b111111111111110010101000100, 27'b111111111111110000010100001, 27'b000000000000001110010110000, 27'b000000000000000100110101100, 27'b111111111111111100000111100, 27'b111111111111110111001111011, 27'b000000000000000101100001000, 27'b000000000000000000000000111, 27'b111111111111111000011001001, 27'b000000000000000000110110011, 27'b000000000000000010001110011, 27'b111111111111111101001010111, 27'b000000000000001001000101101, 27'b111111111111100000101001100, 27'b000000000000000001010011111, 27'b000000000000000111101001100, 27'b111111111111111110101011101, 27'b000000000000000000011110100, 27'b111111111111111000100010010, 27'b111111111111111111111111101, 27'b111111111111111001100100000, 27'b111111111111111111001110101}, 
{27'b000000000000000110110011011, 27'b000000000000001011000010111, 27'b000000000000010001100111111, 27'b111111111111111001011101001, 27'b000000000000001101010100001, 27'b000000000000001001110011010, 27'b000000000000000000000001000, 27'b000000000000001110100100110, 27'b000000000000001011011011011, 27'b111111111111111100100101001, 27'b000000000000010110011100111, 27'b111111111111110100110100110, 27'b000000000000010011111000100, 27'b000000000000001110010010001, 27'b111111111111011101101010100, 27'b111111111111111111111110000, 27'b000000000000000000000000001, 27'b000000000000000000001011110, 27'b000000000000001000010100010, 27'b111111111111101111111001011, 27'b000000000000000111000101111, 27'b111111111111111001001101111, 27'b111111111111110000010011111, 27'b111111111111111010111110110, 27'b000000000000001010100010100, 27'b111111111111101010111000110, 27'b111111111111110101011100101, 27'b111111111111111110101011101, 27'b111111111111111111111111101, 27'b111111111111101101111100010, 27'b000000000000001100101001111, 27'b000000000000000000000000110}, 
{27'b111111111111111110011011000, 27'b000000000000000000000001011, 27'b111111111111111111111111111, 27'b111111111111111111111111111, 27'b111111111111110100110000110, 27'b000000000000000000010010110, 27'b000000000000000000010000111, 27'b111111111111111111100001001, 27'b111111111111111111001110011, 27'b111111111111111110100001110, 27'b000000000000000100011100101, 27'b111111111111111111111110011, 27'b000000000000000010101001110, 27'b111111111111110101000011001, 27'b000000000000000011011010111, 27'b111111111111111111111110100, 27'b000000000000000100100000001, 27'b000000000000001110010100110, 27'b111111111111110100101101101, 27'b000000000000000001101010010, 27'b111111111111111100110101000, 27'b000000000000000100000111011, 27'b000000000000000110000101011, 27'b111111111111111101010001011, 27'b111111111111110111111101100, 27'b000000000000000000101010001, 27'b000000000000011010100010011, 27'b111111111111111111001110011, 27'b111111111111111111100000101, 27'b000000000000001010011000001, 27'b000000000000000000000000011, 27'b000000000000011011100101011}, 
{27'b111111111111101111010011110, 27'b000000000000000001001010000, 27'b111111111111111001000100111, 27'b000000000000001100010000001, 27'b000000000000000011100000101, 27'b111111111111111110111111010, 27'b111111111111111111111111111, 27'b111111111111111111111111111, 27'b111111111111110110010011001, 27'b111111111111111110111100011, 27'b000000000000000000000000010, 27'b111111111111101110001110110, 27'b000000000000000000011001101, 27'b111111111111111110101110100, 27'b111111111111111111111010111, 27'b111111111111111111111111100, 27'b111111111111111100010001000, 27'b000000000000000000001011001, 27'b000000000000000000000110011, 27'b000000000000000101000100111, 27'b000000000000000000100011111, 27'b000000000000000000000000000, 27'b000000000000000000000000010, 27'b111111111111111111101111011, 27'b000000000000000000000000100, 27'b000000000000000000100101100, 27'b000000000000010010100110100, 27'b111111111111111111111111111, 27'b111111111111111111111111101, 27'b111111111111111110101100100, 27'b000000000000000101100110100, 27'b111111111111111111001011110}, 
{27'b111111111111111111111100110, 27'b111111111111111011001010000, 27'b000000000000000110100010011, 27'b000000000000000001010001110, 27'b111111111111110100000110101, 27'b000000000000000000000001001, 27'b000000000000001001001001101, 27'b111111111111111111111111101, 27'b000000000000000000000000000, 27'b111111111111111100110110000, 27'b000000000000000011101011011, 27'b000000000000000000100110111, 27'b000000000000001010010110101, 27'b111111111111101110011101001, 27'b111111111111111100111110011, 27'b111111111111111111011100110, 27'b000000000000000110111010101, 27'b111111111111110011101101011, 27'b000000000000000000101011100, 27'b111111111111100111110110100, 27'b111111111111111111011001010, 27'b111111111111111100001100011, 27'b111111111111111110101101011, 27'b000000000000001001011101100, 27'b111111111111111101100111011, 27'b111111111111110111000000011, 27'b000000000000000010111001000, 27'b000000000000000000000000101, 27'b000000000000001100101010101, 27'b000000000000010000101111100, 27'b111111111111110101100000001, 27'b111111111111110001101000000}, 
{27'b000000000000000010001010001, 27'b000000000000000000110100010, 27'b111111111111110010101111111, 27'b111111111111111110001011110, 27'b111111111111111111111111110, 27'b000000000000000000000100011, 27'b000000000000000011011001101, 27'b000000000000001101001010011, 27'b000000000000000000000000001, 27'b000000000000000000101001100, 27'b000000000000000010001111011, 27'b111111111111101110101111010, 27'b111111111111111101110111101, 27'b111111111111101100101011100, 27'b000000000000001111011000110, 27'b000000000000000000000000110, 27'b111111111111111111111110011, 27'b111111111111101011011111101, 27'b111111111111111111111111011, 27'b111111111111111101100111101, 27'b111111111111111111010101011, 27'b000000000000000000000000000, 27'b000000000000000001111111101, 27'b111111111111111011001100001, 27'b000000000000000001101100110, 27'b000000000000001101001001100, 27'b000000000000001101101001010, 27'b000000000000001100011111111, 27'b000000000000001001110110110, 27'b000000000000000000000000011, 27'b000000000000000011101001111, 27'b000000000000011001000100101}, 
{27'b111111111111111111001100010, 27'b111111111111111000011000111, 27'b000000000000001100011101011, 27'b111111111111111100101101010, 27'b000000000000000010001110111, 27'b000000000000000101010111110, 27'b111111111111111111111111111, 27'b111111111111110110110100010, 27'b111111111111111101010001100, 27'b111111111111101100110001101, 27'b000000000000001110010100000, 27'b000000000000000000000111110, 27'b000000000000001101011010010, 27'b000000000000010101011100011, 27'b111111111111111100010001100, 27'b111111111111100100001000111, 27'b111111111111111100101011010, 27'b000000000000001111000010010, 27'b111111111111110110111100101, 27'b111111111111111001010100101, 27'b000000000000000001111001101, 27'b000000000000000000000010000, 27'b111111111111101110100011110, 27'b111111111111111001111000010, 27'b111111111111111110101111100, 27'b111111111111111100000110100, 27'b000000000000000011100101111, 27'b000000000000010110100000111, 27'b000000000000000111110110110, 27'b111111111111111111111111110, 27'b000000000000000010100101010, 27'b000000000000000000111000100}, 
{27'b000000000000000001010110111, 27'b000000000000001110100001001, 27'b000000000000000000000000001, 27'b000000000000001001011101001, 27'b000000000000011010100110011, 27'b111111111111111010100010010, 27'b111111111111111111111111110, 27'b111111111111111110100101010, 27'b000000000000001001011000000, 27'b111111111111111001110111110, 27'b111111111111111111111101010, 27'b000000000000001010101010101, 27'b000000000000000000010001011, 27'b000000000000000000111000001, 27'b111111111111001111001000101, 27'b111111111111111101011101011, 27'b000000000000000000000000000, 27'b000000000000000110011011000, 27'b111111111111111111111001001, 27'b000000000000001001100011100, 27'b111111111111111111111111100, 27'b111111111111111010011110001, 27'b111111111111101110000001001, 27'b000000000000000100001011111, 27'b000000000000001001001001100, 27'b111111111111011100100000011, 27'b111111111111111111111111100, 27'b000000000000000000000000010, 27'b000000000000010001011010010, 27'b111111111111100110010110110, 27'b000000000000000000000011101, 27'b111111111111111111110011100}, 
{27'b000000000000000000010011010, 27'b111111111111110101001000011, 27'b000000000000000001101110100, 27'b111111111111111111100001011, 27'b000000000000000001101010101, 27'b000000000000010000111011100, 27'b111111111111101000110011101, 27'b000000000000000001000110011, 27'b000000000000001101100011001, 27'b111111111111110101001101011, 27'b111111111111111111010000011, 27'b000000000000000001100100001, 27'b111111111111111111101101101, 27'b000000000000000101101110010, 27'b000000000000000011011011111, 27'b111111111111111111011101111, 27'b000000000000000010001001010, 27'b000000000000000000000000100, 27'b000000000000000000101100001, 27'b000000000000001100001001111, 27'b111111111111111111000110100, 27'b111111111111110000100000000, 27'b111111111111101100101001001, 27'b111111111111111001110011010, 27'b111111111111101101000110010, 27'b000000000000000110101010000, 27'b000000000000010011111100011, 27'b000000000000001011110011000, 27'b111111111111111111101010101, 27'b111111111111110100000100111, 27'b111111111111110110000011100, 27'b000000000000000001111010010}, 
{27'b000000000000000001101010010, 27'b111111111111110000101101110, 27'b111111111111111111011101011, 27'b000000000000000100110100001, 27'b111111111111110000101100000, 27'b000000000000000101011011100, 27'b111111111111111111111111110, 27'b111111111111111111111111101, 27'b111111111111111111111111111, 27'b000000000000000000000000011, 27'b000000000000001000011101011, 27'b111111111111111111011100101, 27'b000000000000000000010011111, 27'b000000000000000000000000100, 27'b000000000000000100000100110, 27'b111111111111111111011101011, 27'b000000000000000000000101101, 27'b111111111111111111111110100, 27'b111111111111110101101100011, 27'b111111111111101111110100011, 27'b111111111111111111111110110, 27'b111111111111101110111010101, 27'b111111111111110110010111001, 27'b111111111111110100000110101, 27'b000000000000011100011111111, 27'b000000000000000000100100000, 27'b111111111111111110100001101, 27'b000000000000001010001001111, 27'b000000000000011100101110000, 27'b000000000000001100101000101, 27'b111111111111011110000100001, 27'b111111111111111010000100000}, 
{27'b000000000000001100000001110, 27'b111111111111111111111111001, 27'b000000000000001000000010000, 27'b111111111111111111010111010, 27'b000000000000001111011110101, 27'b111111111111111011011011111, 27'b000000000000000010010001000, 27'b000000000000001101011000100, 27'b000000000000001000100100011, 27'b111111111111101111010010100, 27'b111111111111111110000001111, 27'b000000000000000011111011101, 27'b000000000000000010001101001, 27'b111111111111111111100010000, 27'b000000000000000010101101111, 27'b000000000000000000000000100, 27'b000000000000001011100110001, 27'b000000000000000001000111110, 27'b000000000000001011111110010, 27'b111111111111111101111001110, 27'b111111111111111011111011001, 27'b111111111111111101100110110, 27'b111111111111111111111111100, 27'b000000000000001001101010001, 27'b111111111111111001100001100, 27'b111111111111111111110011010, 27'b000000000000000000000000000, 27'b000000000000000000000000100, 27'b000000000000000000000000010, 27'b000000000000001001010110001, 27'b111111111111110101101111010, 27'b111111111111111111010000011}, 
{27'b111111111111111111111110101, 27'b111111111111111111000000110, 27'b111111111111110001000111100, 27'b000000000000001001000110101, 27'b000000000000000111001001000, 27'b111111111111111100011111100, 27'b111111111111111111111111101, 27'b111111111111111000101111010, 27'b000000000000000000001101110, 27'b111111111111111111111111010, 27'b111111111111110110010110110, 27'b111111111111111000000111100, 27'b000000000000001111010101000, 27'b000000000000000000000000000, 27'b111111111111111011111010011, 27'b111111111111111111111111111, 27'b000000000000000110110110011, 27'b111111111111111111111111101, 27'b111111111111111111111111111, 27'b111111111111111001000101101, 27'b000000000000001010000111110, 27'b000000000000000000000000001, 27'b000000000000000100111111110, 27'b111111111111111111000101010, 27'b000000000000000101000001100, 27'b000000000000000000000100100, 27'b000000000000000000000000001, 27'b000000000000000111101101000, 27'b111111111111111001110110100, 27'b111111111111111110100001101, 27'b000000000000000101001000110, 27'b111111111111111100100111001}, 
{27'b111111111111111111011101101, 27'b111111111111110110001000000, 27'b000000000000010011000001010, 27'b111111111111111101111010111, 27'b000000000000000110010010001, 27'b111111111111110110110110000, 27'b000000000000000000000000001, 27'b000000000000000001000110000, 27'b111111111111110000101010111, 27'b111111111111111111100101110, 27'b111111111111111100000010100, 27'b000000000000000001110111001, 27'b111111111111110101100000011, 27'b000000000000000100011010011, 27'b000000000000000110011110010, 27'b000000000000000011100000011, 27'b000000000000000010101111101, 27'b111111111111111110110010000, 27'b111111111111101001010101101, 27'b111111111111111111100100011, 27'b111111111111111110001011011, 27'b000000000000000100011110011, 27'b111111111111111100011100100, 27'b111111111111111111111111111, 27'b000000000000000110010100111, 27'b111111111111111110100010101, 27'b111111111111111111100010011, 27'b000000000000001100011100101, 27'b111111111111110011010000111, 27'b111111111111110110100011100, 27'b000000000000001011001110011, 27'b000000000000000001001001100}, 
{27'b000000000000001101110010100, 27'b000000000000000110011100010, 27'b000000000000000000000001100, 27'b111111111111111010111010011, 27'b111111111111111101011111010, 27'b111111111111111111111110010, 27'b000000000000000000000000001, 27'b111111111111111101110010011, 27'b111111111111111100000001101, 27'b111111111111111100001101010, 27'b000000000000000000000000101, 27'b000000000000000101000100010, 27'b000000000000000000001101000, 27'b000000000000000001101100010, 27'b111111111111111110100100100, 27'b000000000000000000001011110, 27'b111111111111111011000101111, 27'b000000000000000000000001001, 27'b111111111111111111011011111, 27'b111111111111111111111110110, 27'b000000000000000000000100110, 27'b000000000000000001111001101, 27'b000000000000000011000111000, 27'b000000000000000000000000001, 27'b000000000000000000000000100, 27'b111111111111101100011101101, 27'b111111111111111001100111111, 27'b000000000000000000001101100, 27'b000000000000000000101001111, 27'b000000000000000000000010101, 27'b111111111111111010010101010, 27'b000000000000000000101011111}, 
{27'b000000000000000110000000010, 27'b111111111111011110100100110, 27'b111111111111111111111111110, 27'b111111111111111101100101111, 27'b111111111111111000100011000, 27'b111111111111111111101100010, 27'b000000000000000000000000000, 27'b000000000000010001100001111, 27'b111111111111111110100110010, 27'b111111111111111111010011000, 27'b000000000000000010101000111, 27'b111111111111101010110110111, 27'b000000000000000000110001001, 27'b111111111111110001111110000, 27'b000000000000010111000111100, 27'b111111111111111110010100111, 27'b111111111111111000110000001, 27'b111111111111101110011111101, 27'b111111111111111111101010011, 27'b111111111111101001010110011, 27'b111111111111100110000101110, 27'b111111111111111111111111011, 27'b000000000000000000000000111, 27'b000000000000000000000000001, 27'b000000000000000111110011110, 27'b111111111111111111100011011, 27'b111111111111110110011101010, 27'b111111111111111101101011001, 27'b111111111111111111010000010, 27'b000000000000000000000000011, 27'b111111111111111110111111000, 27'b111111111111101001100110100}
};

localparam logic signed [26:0] bias [32] = '{
27'b000000000000001000011100110,  // 0.5280959606170654
27'b000000000000001101011101101,  // 0.8414360880851746
27'b000000000000000110010111011,  // 0.397830605506897
27'b000000000000000110100100011,  // 0.4105983078479767
27'b111111111111000101011110011,  // -3.657735586166382
27'b111111111111110001101000101,  // -0.8977976441383362
27'b000000000000011011010010000,  // 1.7051936388015747
27'b111111111111101011100100110,  // -1.2765135765075684
27'b111111111111110110101010001,  // -0.5837795734405518
27'b000000000000101011001100011,  // 2.699671983718872
27'b000000000000000011011110010,  // 0.2170683741569519
27'b000000000000001110000110100,  // 0.8814588785171509
27'b111111111111010101110110011,  // -2.634300947189331
27'b111111111111100001111101101,  // -1.877297282218933
27'b000000000000011010100110011,  // 1.6625694036483765
27'b000000000000101011111011110,  // 2.7459704875946045
27'b111111111111111000010110001,  // -0.47838035225868225
27'b000000000000011011001011010,  // 1.6984987258911133
27'b000000000000001101101011011,  // 0.8548859357833862
27'b000000000000010000000100101,  // 1.0045719146728516
27'b000000000000010110101101110,  // 1.4197649955749512
27'b000000000000001101010100011,  // 0.832463800907135
27'b000000000000001000101100011,  // 0.5434179306030273
27'b000000000000001110110101111,  // 0.9277304410934448
27'b111111111111111010100001001,  // -0.3426123857498169
27'b111111111111110111000011111,  // -0.5587119460105896
27'b111111111111110110000100001,  // -0.6208624839782715
27'b111111111111101011100001000,  // -1.2802538871765137
27'b000000000000000000111100110,  // 0.05940237268805504
27'b111111111111110010110110111,  // -0.8213341236114502
27'b000000000000001110000011011,  // 0.8783953189849854
27'b111111111111110000110011100   // -0.949700653553009
};
endpackage