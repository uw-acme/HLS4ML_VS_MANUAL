// Width: 21
// NFRAC: 10
package dense_1_21_10;

localparam logic signed [20:0] weights [16][64] = '{ 
{21'b000000000000100000101, 21'b111111111110101100100, 21'b111111111111101000110, 21'b111111111111100011000, 21'b111111111111001100001, 21'b000000000000001110001, 21'b111111111101111011010, 21'b000000000000000000000, 21'b000000000000000111011, 21'b000000000000100001101, 21'b000000000000000000011, 21'b111111111111001100001, 21'b111111111111111111110, 21'b000000000000011010110, 21'b000000000000000100010, 21'b111111111111011110100, 21'b000000000000011101110, 21'b000000000000000111100, 21'b000000000000000000000, 21'b111111111111111111111, 21'b000000000000110000001, 21'b111111111111010101100, 21'b111111111111111101001, 21'b000000000000111100100, 21'b111111111111010110110, 21'b111111111110101000101, 21'b111111111111011100101, 21'b111111111111100111000, 21'b111111111111110010100, 21'b111111111111111111110, 21'b000000000000000100110, 21'b000000000000011111011, 21'b000000000000011001000, 21'b111111111111111110010, 21'b000000000000000000000, 21'b000000000000100111110, 21'b111111111111111101101, 21'b111111111111011111110, 21'b000000000000000011011, 21'b000000000000011000101, 21'b111111111111111110011, 21'b000000000000100011001, 21'b111111111111011101111, 21'b000000000001110110111, 21'b111111111111111111110, 21'b000000000000111001111, 21'b000000000000000000000, 21'b000000000000010111100, 21'b000000000000011001000, 21'b111111111111111100111, 21'b000000000000000000000, 21'b000000000000010100100, 21'b000000000000011011101, 21'b000000000000001001111, 21'b111111111111110001001, 21'b111111111111011000010, 21'b000000000001000100101, 21'b111111111111000000000, 21'b000000000000111011110, 21'b111111111111010010101, 21'b000000000001100101100, 21'b111111111111111111000, 21'b000000000000000001011, 21'b000000000000001010011}, 
{21'b000000000000000000010, 21'b111111111111010110111, 21'b111111111111101111000, 21'b111111111111011100001, 21'b111111111111010111010, 21'b000000000000001101101, 21'b111111111110011111011, 21'b111111111111111111101, 21'b111111111111100010111, 21'b000000000000010110000, 21'b000000000000000000110, 21'b111111111111110100111, 21'b000000000000011001001, 21'b000000000000000000000, 21'b111111111111111111111, 21'b000000000000011010100, 21'b111111111111111111001, 21'b000000000000000000000, 21'b111111111111101000101, 21'b111111111111011111111, 21'b000000000000111000100, 21'b111111111111110101101, 21'b000000000000000110001, 21'b000000000001011001011, 21'b000000000000100000111, 21'b111111111111100010100, 21'b111111111111100010011, 21'b111111111111111111111, 21'b111111111111110011000, 21'b111111111111001100000, 21'b111111111111111000010, 21'b000000000000111010001, 21'b000000000000100011101, 21'b000000000001000110011, 21'b000000000001010000100, 21'b000000000000000110011, 21'b111111111111110000110, 21'b111111111111001000011, 21'b000000000000000111010, 21'b000000000000011000001, 21'b000000000000000010111, 21'b000000000000011010011, 21'b111111111111100100110, 21'b000000000000100000010, 21'b000000000000010110000, 21'b000000000000000110011, 21'b111111111111010100011, 21'b000000000000001010001, 21'b000000000000100001010, 21'b000000000000000011110, 21'b000000000000000011001, 21'b000000000010010100001, 21'b111111111111110110011, 21'b111111111111110011011, 21'b111111111111111001000, 21'b111111111111111111000, 21'b000000000000100000111, 21'b111111111111010000101, 21'b000000000001111110000, 21'b000000000000000000100, 21'b000000000001000010101, 21'b000000000000011110101, 21'b000000000001101001010, 21'b000000000000010010000}, 
{21'b111111111111111111000, 21'b000000000000000000000, 21'b111111111111110101010, 21'b111111111111101001011, 21'b111111111111101000010, 21'b000000000000000101010, 21'b000000000010111101100, 21'b111111111111111111111, 21'b111111111101011101111, 21'b111111111111111111111, 21'b111111111111111111110, 21'b111111111111111101101, 21'b111111111111100010111, 21'b000000000000000000001, 21'b111111111111111110110, 21'b000000000000010101100, 21'b000000000001110011111, 21'b111111111111111111111, 21'b000000000000001001001, 21'b000000000000000000000, 21'b000000000000110100110, 21'b111111111110100011101, 21'b000000000001001001111, 21'b111111111110100100101, 21'b000000000001111001011, 21'b111111111111010011101, 21'b111111111111100000101, 21'b111111111110100100001, 21'b000000000010100011000, 21'b000000000000100011010, 21'b000000000000000001011, 21'b000000000001000010010, 21'b000000000010000010100, 21'b111111111101100111000, 21'b111111111111110011110, 21'b000000000000000100000, 21'b111111111111100010011, 21'b000000000001110010110, 21'b111111111111111010111, 21'b000000000000101000000, 21'b000000000000101010101, 21'b000000000000101111010, 21'b111111111111111111111, 21'b111111111111111111111, 21'b111111111111111101110, 21'b000000000000010100000, 21'b111111111111011100001, 21'b111111111111101010001, 21'b111111111111111101110, 21'b000000000000110010010, 21'b111111111111101001011, 21'b000000000000010011001, 21'b111111111111111111111, 21'b000000000000010001001, 21'b111111111111101001100, 21'b111111111111111111111, 21'b111111111111011000100, 21'b111111111110101010010, 21'b111111111111111111101, 21'b000000000000000000000, 21'b000000000011000101011, 21'b000000000000000001101, 21'b111111111111111111101, 21'b111111111111011000011}, 
{21'b111111111111000101010, 21'b111111111111010000110, 21'b111111111110100111010, 21'b000000000000100111011, 21'b111111111111010111100, 21'b111111111101010011101, 21'b111111111111110001010, 21'b111111111111011000100, 21'b000000000000011100101, 21'b111111111111111111111, 21'b000000000010100001111, 21'b111111111111110010011, 21'b111111111110011011110, 21'b000000000001001010001, 21'b000000000000000011001, 21'b111111111111111111110, 21'b111111111111000111001, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111100011000, 21'b111111111101101100101, 21'b111111111111110001101, 21'b111111111110100110100, 21'b000000000000011001011, 21'b111111111111001110011, 21'b111111111110001010001, 21'b000000000000101000000, 21'b000000000001011110010, 21'b000000000010100101110, 21'b111111111111000101001, 21'b111111111110110101011, 21'b000000000000001001011, 21'b000000000001000000000, 21'b111111111110010100010, 21'b111111111111010111110, 21'b000000000000000000000, 21'b111111111110100011000, 21'b000000000000011111000, 21'b111111111111000111100, 21'b000000000000001111010, 21'b000000000000111010101, 21'b000000000000010100000, 21'b000000000000000000000, 21'b000000000000000010100, 21'b000000000001000110101, 21'b111111111111100110011, 21'b111111111111111111111, 21'b111111111111010011111, 21'b111111111111111111111, 21'b111111111111110011100, 21'b111111111110110001001, 21'b000000000000001011000, 21'b111111111111111111111, 21'b000000000000011011111, 21'b000000000000101000010, 21'b000000000001010010110, 21'b111111111110000100001, 21'b111111111110001001000, 21'b111111111110100101101, 21'b000000000001101110111, 21'b000000000011011111111, 21'b111111111110001100110, 21'b111111111111111001000, 21'b000000000000110111100}, 
{21'b000000000000101011110, 21'b111111111110110000110, 21'b111111111111011110110, 21'b111111111111111111111, 21'b111111111111101100010, 21'b000000000000101011100, 21'b000000000000011000010, 21'b111111111111111111111, 21'b111111111110110011100, 21'b111111111111100001000, 21'b111111111111010000110, 21'b000000000000000110110, 21'b000000000000000000001, 21'b000000000000000000000, 21'b111111111111111010110, 21'b000000000000101101110, 21'b000000000000010001000, 21'b111111111111001101101, 21'b000000000000000011111, 21'b000000000000000001101, 21'b000000000000011010111, 21'b111111111111110000111, 21'b000000000000001001100, 21'b111111111111111101100, 21'b000000000010001000011, 21'b111111111111101000001, 21'b111111111111011100000, 21'b111111111111001100010, 21'b000000000000000000000, 21'b000000000000010101000, 21'b000000000000001110111, 21'b000000000000100011000, 21'b111111111111111110011, 21'b000000000000001001011, 21'b000000000000010000101, 21'b111111111111111111111, 21'b000000000000000000110, 21'b000000000001110000110, 21'b111111111111011011000, 21'b111111111111110110001, 21'b000000000000110111011, 21'b000000000000011111110, 21'b111111111111000001011, 21'b000000000000000000110, 21'b111111111101110111010, 21'b111111111111111111111, 21'b111111111111110000010, 21'b000000000000000001100, 21'b111111111111111111111, 21'b111111111111111100111, 21'b111111111111111111111, 21'b000000000000011000000, 21'b111111111111111111010, 21'b000000000000101000101, 21'b111111111111100111100, 21'b111111111110100001111, 21'b111111111111000100010, 21'b111111111110111110110, 21'b111111111110110001011, 21'b000000000001011111100, 21'b000000000010101111110, 21'b000000000001100101011, 21'b000000000000001111101, 21'b111111111111111111111}, 
{21'b111111111111000110111, 21'b111111111110101111010, 21'b000000000000000000000, 21'b000000000000100111010, 21'b000000000000100100100, 21'b111111111111100100110, 21'b000000000001001010100, 21'b111111111111111111111, 21'b000000000000011111001, 21'b111111111111111111111, 21'b111111111111111110110, 21'b111111111111110110101, 21'b111111111111101001011, 21'b000000000001001010000, 21'b111111111111110100100, 21'b000000000000000000000, 21'b111111111110110000000, 21'b111111111111010010101, 21'b000000000000000000000, 21'b111111111111111111111, 21'b111111111111111001111, 21'b111111111111010111110, 21'b111111111111010111001, 21'b000000000000111011100, 21'b111111111111010111010, 21'b111111111111111111111, 21'b000000000000100000110, 21'b111111111111110110101, 21'b111111111110001000100, 21'b111111111111111111111, 21'b111111111111110111011, 21'b111111111111111110101, 21'b111111111111111110100, 21'b000000000000000101001, 21'b000000000000010000111, 21'b000000000000101100010, 21'b000000000000000001101, 21'b111111111111110011011, 21'b111111111111011110011, 21'b111111111111111111110, 21'b111111111111101010010, 21'b111111111110111100111, 21'b000000000000110011001, 21'b000000000000000001011, 21'b000000000001001101001, 21'b000000000000000000000, 21'b111111111111111111111, 21'b000000000000001100001, 21'b111111111111001010010, 21'b000000000000011101111, 21'b000000000000000000000, 21'b111111111111110011000, 21'b111111111111010001101, 21'b000000000000110001011, 21'b111111111111111111111, 21'b000000000000101100011, 21'b000000000000011011101, 21'b000000000000011010000, 21'b111111111111111101100, 21'b111111111111111110111, 21'b111111111110011000100, 21'b111111111111101111110, 21'b111111111111111000101, 21'b111111111111111111111}, 
{21'b111111111111011011110, 21'b111111111111010101000, 21'b111111111111001000110, 21'b111111111111110111000, 21'b111111111111101110111, 21'b000000000000001101010, 21'b111111111110100110101, 21'b111111111111101100110, 21'b111111111111100011010, 21'b111111111111111111111, 21'b111111111111011011001, 21'b000000000000101100100, 21'b000000000000000100100, 21'b000000000000010001101, 21'b000000000000100111111, 21'b000000000000000000000, 21'b000000000001100110000, 21'b000000000000001011011, 21'b000000000000011111000, 21'b000000000000100010010, 21'b111111111111101011111, 21'b000000000000101110100, 21'b111111111111100000111, 21'b111111111110111111110, 21'b000000000000010110001, 21'b000000000001000010001, 21'b111111111111111111011, 21'b000000000000000110111, 21'b111111111110000110010, 21'b000000000000100100101, 21'b000000000000100010001, 21'b111111111111010000001, 21'b000000000000111100010, 21'b000000000001010101000, 21'b000000000000000000000, 21'b000000000000101011110, 21'b111111111111111111111, 21'b000000000000100100011, 21'b000000000000011001011, 21'b000000000000000000000, 21'b111111111111110000111, 21'b111111111111010001011, 21'b000000000000010010010, 21'b000000000000111101110, 21'b000000000001000010011, 21'b111111111111101010011, 21'b111111111111110101010, 21'b111111111111100111101, 21'b111111111111101110101, 21'b000000000000001111001, 21'b000000000000000000011, 21'b000000000000000100010, 21'b000000000000000000000, 21'b000000000000010111001, 21'b111111111111101001101, 21'b000000000001100010101, 21'b000000000000101101100, 21'b111111111111111100110, 21'b000000000000110001111, 21'b000000000000011011110, 21'b111111111100101111111, 21'b111111111110110110001, 21'b111111111111101001111, 21'b111111111111111110101}, 
{21'b000000000000000000101, 21'b000000000000011110100, 21'b111111111111111111111, 21'b111111111111111111111, 21'b111111111111010110110, 21'b111111111111111100000, 21'b111111111111011111000, 21'b000000000000000000000, 21'b000000000000000011100, 21'b000000000000110001110, 21'b000000000000000001110, 21'b111111111111001111101, 21'b111111111111110111111, 21'b000000000000000000000, 21'b111111111111111001010, 21'b111111111111000110011, 21'b111111111110010011011, 21'b111111111111111111111, 21'b111111111110110010101, 21'b111111111111000110111, 21'b111111111111001110001, 21'b000000000000101100011, 21'b000000000000000110000, 21'b111111111111101101110, 21'b111111111111001000000, 21'b000000000000010011111, 21'b000000000000000000000, 21'b000000000000111111111, 21'b000000000001100111001, 21'b111111111111111010110, 21'b000000000000000000000, 21'b000000000000011101100, 21'b111111111110101000101, 21'b111111111111010000100, 21'b000000000000000111000, 21'b000000000000001011110, 21'b111111111111011100000, 21'b000000000000011110101, 21'b000000000000010000111, 21'b111111111111101100011, 21'b111111111111001010010, 21'b111111111111111011010, 21'b000000000000000100001, 21'b111111111111101010101, 21'b000000000000000111001, 21'b000000000000011101010, 21'b111111111111110000101, 21'b000000000000000011000, 21'b000000000000000000000, 21'b111111111111100100000, 21'b111111111111001110010, 21'b000000000000110101001, 21'b000000000000010000001, 21'b111111111111101001001, 21'b000000000000010000111, 21'b111111111111111000000, 21'b111111111111000011010, 21'b111111111111101110111, 21'b111111111111111001010, 21'b111111111111110111000, 21'b000000000001101010010, 21'b000000000000011000011, 21'b111111111111111001110, 21'b111111111111111111111}, 
{21'b000000000000000001111, 21'b000000000001001011000, 21'b111111111110110101101, 21'b111111111111100010011, 21'b000000000000101001010, 21'b111111111111100101100, 21'b000000000010011011000, 21'b111111111111011011001, 21'b111111111111111111111, 21'b000000000000100101100, 21'b000000000000100000100, 21'b111111111111111111101, 21'b111111111111111001110, 21'b111111111111000010010, 21'b000000000000100100000, 21'b000000000000010100011, 21'b111111111111100111001, 21'b111111111111111111111, 21'b000000000000000000000, 21'b000000000000000000000, 21'b000000000000100001111, 21'b111111111111000101001, 21'b000000000000110010001, 21'b000000000001001110011, 21'b111111111111110100110, 21'b111111111111111111111, 21'b111111111111111101111, 21'b111111111111111111111, 21'b000000000001011110001, 21'b000000000000000000101, 21'b111111111111011101000, 21'b000000000000000000000, 21'b000000000000110001001, 21'b111111111110011000001, 21'b111111111110111010110, 21'b000000000000011001011, 21'b000000000000010001101, 21'b111111111110110110110, 21'b111111111111100111110, 21'b111111111111100100100, 21'b000000000000110011010, 21'b000000000000110010000, 21'b000000000000000000000, 21'b111111111111011101011, 21'b000000000000000000000, 21'b000000000000110010100, 21'b111111111111111000011, 21'b111111111111111111111, 21'b000000000000000001011, 21'b000000000000011111010, 21'b111111111111111000101, 21'b111111111111100111001, 21'b000000000000101100000, 21'b111111111111100100011, 21'b000000000000100011110, 21'b000000000001001010110, 21'b000000000000000101000, 21'b000000000000100001101, 21'b111111111111001100110, 21'b111111111111010001000, 21'b000000000001101010011, 21'b111111111111101111100, 21'b000000000000000101111, 21'b111111111111110100000}, 
{21'b000000000000000010000, 21'b111111111111000110000, 21'b000000000000101111001, 21'b111111111111011011101, 21'b111111111111111111100, 21'b000000000000011011000, 21'b111111111110110101100, 21'b000000000000011000100, 21'b000000000000111110110, 21'b000000000000010011101, 21'b000000000000101110011, 21'b000000000000101001010, 21'b111111111111011000111, 21'b111111111111110110010, 21'b111111111111111001011, 21'b000000000000000000001, 21'b111111111110000101001, 21'b000000000000101001010, 21'b111111111111111011010, 21'b000000000000000011111, 21'b111111111111010010111, 21'b000000000000001000111, 21'b000000000000010011100, 21'b111111111111111111111, 21'b111111111111000101000, 21'b111111111111111001111, 21'b111111111111110101100, 21'b000000000010011111101, 21'b111111111110101011001, 21'b000000000000001000100, 21'b000000000000001100011, 21'b111111111111111000100, 21'b111111111111100011101, 21'b000000000000001110111, 21'b111111111111110101111, 21'b111111111111101110110, 21'b111111111111101001001, 21'b111111111111100101000, 21'b111111111111111101001, 21'b111111111111011001111, 21'b000000000000101001001, 21'b000000000000001111110, 21'b000000000000111111100, 21'b000000000000001011001, 21'b000000000000000100101, 21'b111111111111011010110, 21'b000000000000000000000, 21'b111111111111111111111, 21'b111111111111111111111, 21'b000000000000011000110, 21'b000000000000010110101, 21'b000000000000100101101, 21'b111111111111111111001, 21'b111111111111011010011, 21'b000000000000000001001, 21'b000000000000000000000, 21'b000000000000101001010, 21'b111111111111100110010, 21'b111111111110111001100, 21'b000000000001000111110, 21'b111111111111011010011, 21'b000000000010010100111, 21'b111111111111111101011, 21'b111111111111010010101}, 
{21'b111111111110110110001, 21'b111111111111111111110, 21'b111111111111001011100, 21'b000000000000011101011, 21'b000000000000100001101, 21'b111111111111110010111, 21'b000000000001000010001, 21'b111111111111101010001, 21'b111111111111000010101, 21'b111111111111010001000, 21'b111111111111011111110, 21'b111111111111000011000, 21'b111111111111100010101, 21'b000000000000011001001, 21'b000000000000000000000, 21'b000000000000000000000, 21'b000000000001101011110, 21'b111111111111111010011, 21'b111111111111111111110, 21'b000000000000110100101, 21'b000000000000100101011, 21'b111111111110110101111, 21'b111111111111001111000, 21'b000000000000011000001, 21'b111111111111001000111, 21'b111111111111111101010, 21'b111111111111011110110, 21'b111111111111010101001, 21'b111111111111001000001, 21'b000000000000100110101, 21'b000000000000011101001, 21'b111111111111101100000, 21'b111111111111110110101, 21'b111111111110000011010, 21'b111111111111101001011, 21'b000000000000000110010, 21'b111111111111101111011, 21'b111111111111011010000, 21'b111111111111111111100, 21'b000000000000001111001, 21'b111111111111110000110, 21'b111111111111111111101, 21'b111111111111111011100, 21'b111111111110101010111, 21'b000000000000000000000, 21'b000000000000000000000, 21'b000000000000101011100, 21'b111111111111110000000, 21'b000000000000110110001, 21'b111111111111100111100, 21'b000000000000100100110, 21'b111111111111111111110, 21'b000000000000011100111, 21'b111111111111001101111, 21'b111111111111111111111, 21'b000000000001000001100, 21'b000000000000101000000, 21'b000000000000100101011, 21'b000000000000000011001, 21'b111111111111001100110, 21'b111111111111011001101, 21'b111111111110101000001, 21'b111111111111111111110, 21'b000000000000001101101}, 
{21'b000000000000100111011, 21'b000000000000000000010, 21'b000000000000010000110, 21'b111111111111111111111, 21'b000000000000010011101, 21'b111111111111101110110, 21'b000000000000011110000, 21'b000000000000000101011, 21'b000000000000010001011, 21'b000000000000101011100, 21'b111111111111011110010, 21'b111111111111111101010, 21'b111111111111111110111, 21'b111111111111111110111, 21'b111111111110101011100, 21'b111111111111011001111, 21'b000000000001010000101, 21'b111111111111111100011, 21'b111111111111111001010, 21'b000000000000000000000, 21'b111111111111001111010, 21'b000000000000000001001, 21'b000000000000100000000, 21'b000000000000000100110, 21'b000000000000000100101, 21'b000000000000101011010, 21'b000000000000000000000, 21'b000000000000000100110, 21'b000000000000000000000, 21'b111111111111111001111, 21'b111111111111100110010, 21'b111111111110101010110, 21'b000000000000100001110, 21'b000000000000101011111, 21'b111111111111111100010, 21'b111111111111100001111, 21'b000000000000000000000, 21'b111111111110101100001, 21'b111111111111111010001, 21'b111111111111111111100, 21'b000000000000011001000, 21'b111111111111101111010, 21'b111111111111111111111, 21'b000000000001101100011, 21'b000000000000111001011, 21'b111111111111111111001, 21'b111111111111111111111, 21'b111111111111111111111, 21'b111111111111100001001, 21'b000000000000010010110, 21'b000000000000010010011, 21'b000000000000010110010, 21'b000000000000010100001, 21'b000000000000110001101, 21'b000000000000101100110, 21'b000000000001010100011, 21'b111111111111101110000, 21'b000000000000110010010, 21'b000000000000010011100, 21'b111111111111010110010, 21'b000000000000001110001, 21'b111111111111001110010, 21'b111111111111000111101, 21'b111111111111000000001}, 
{21'b000000000000000000000, 21'b000000000000011101001, 21'b111111111111100111000, 21'b000000000000000000000, 21'b111111111111111001101, 21'b111111111111111011101, 21'b111111111110101011011, 21'b111111111111111111111, 21'b000000000000100000011, 21'b000000000000011111111, 21'b000000000000011110011, 21'b111111111111001101000, 21'b111111111111110100100, 21'b000000000000100100010, 21'b111111111111111111111, 21'b000000000000000000100, 21'b111111111110010100010, 21'b111111111111111111111, 21'b000000000000101111101, 21'b000000000000001001000, 21'b000000000000011110011, 21'b111111111111110001001, 21'b000000000000011111111, 21'b000000000000110011110, 21'b111111111111010010100, 21'b111111111111011100001, 21'b111111111111111111010, 21'b111111111111110101101, 21'b000000000000001000100, 21'b000000000000000000000, 21'b111111111111111111111, 21'b000000000000101000001, 21'b111111111110100000000, 21'b000000000000101110010, 21'b000000000001000000001, 21'b000000000000001110111, 21'b000000000000001110011, 21'b111111111111110010001, 21'b000000000000001110101, 21'b111111111111110010010, 21'b111111111111011111110, 21'b111111111111111001100, 21'b000000000000010101000, 21'b000000000001011001100, 21'b111111111110010011100, 21'b111111111111000110111, 21'b000000000000011000100, 21'b111111111111110011011, 21'b000000000000111001101, 21'b111111111111100001110, 21'b111111111111010101101, 21'b111111111111011100001, 21'b111111111111111111111, 21'b000000000000001111011, 21'b111111111111101011110, 21'b111111111110010100111, 21'b111111111111101101101, 21'b111111111111111110101, 21'b000000000000000101100, 21'b111111111110110001111, 21'b000000000010001111010, 21'b111111111110111010010, 21'b000000000001000101010, 21'b000000000000010011100}, 
{21'b000000000000001010000, 21'b111111111111100111011, 21'b000000000001010000011, 21'b111111111111011001010, 21'b111111111111000100101, 21'b000000000000001011100, 21'b000000000000100111100, 21'b000000000000100110011, 21'b111111111111101001010, 21'b111111111111101011011, 21'b000000000000000110101, 21'b000000000000011101010, 21'b000000000000011110000, 21'b000000000000000110011, 21'b111111111111100101110, 21'b000000000000010000011, 21'b000000000000111100010, 21'b111111111111111110100, 21'b111111111111011100001, 21'b000000000000000000000, 21'b000000000000001001100, 21'b000000000000000010100, 21'b111111111111011010011, 21'b000000000000001110011, 21'b000000000001100100101, 21'b000000000000000001010, 21'b000000000000010111000, 21'b111111111110011010011, 21'b111111111111110110101, 21'b000000000000000001001, 21'b111111111111100110111, 21'b111111111111011000000, 21'b000000000000111010101, 21'b111111111111111100100, 21'b111111111111111011001, 21'b111111111111011000111, 21'b000000000000010001101, 21'b000000000000100101011, 21'b111111111111111110110, 21'b111111111111111010011, 21'b111111111111101000000, 21'b000000000000011101001, 21'b000000000000000000000, 21'b111111111110101000001, 21'b000000000000100111110, 21'b000000000000110011000, 21'b111111111111111111111, 21'b000000000000000011010, 21'b111111111111001000011, 21'b111111111111110110011, 21'b111111111111111111111, 21'b111111111111010111010, 21'b000000000000000000000, 21'b111111111111101001111, 21'b000000000000000111010, 21'b111111111110010111011, 21'b111111111111111111111, 21'b111111111111111111111, 21'b000000000000100011001, 21'b000000000001001000000, 21'b111111111110100111000, 21'b000000000001000010100, 21'b000000000000000100101, 21'b111111111111110110011}, 
{21'b000000000000100100110, 21'b000000000010011110110, 21'b000000000000111111011, 21'b000000000000100100100, 21'b111111111111000010110, 21'b111111111111010111010, 21'b111111111010110011010, 21'b111111111111000101100, 21'b000000000000110011100, 21'b111111111111111111111, 21'b000000000000100101101, 21'b000000000001101110011, 21'b000000000000001000111, 21'b000000000000000000101, 21'b111111111111111101110, 21'b000000000000000000000, 21'b111111111111100111110, 21'b111111111111100110000, 21'b000000000000011101011, 21'b111111111110111111101, 21'b111111111110101010111, 21'b111111111111110010110, 21'b111111111110110101010, 21'b000000000000000011110, 21'b111111111011011100100, 21'b000000000001101000010, 21'b000000000001111110100, 21'b000000000001001101010, 21'b111111111100100000110, 21'b111111111111010111111, 21'b111111111110100111111, 21'b111111111110010100000, 21'b111111111010111100110, 21'b000000000001010110100, 21'b111111111111111010011, 21'b000000000000101000110, 21'b000000000000000011000, 21'b111111111101001000100, 21'b000000000000000000000, 21'b000000000000000000000, 21'b000000000000000100000, 21'b000000000010000010011, 21'b111111111111100101110, 21'b111111111110101101011, 21'b000000000001110010110, 21'b111111111111000111001, 21'b111111111111010110011, 21'b111111111111001101110, 21'b000000000000111101000, 21'b000000000001000100000, 21'b111111111111110111010, 21'b111111111111010011010, 21'b111111111111111111101, 21'b111111111111110001100, 21'b000000000000000000000, 21'b111111111111001111101, 21'b000000000001001101101, 21'b000000000010001010110, 21'b000000000001011011000, 21'b111111111110001011101, 21'b111111111000100110000, 21'b000000000001110001010, 21'b000000000000001011110, 21'b000000000000101000100}, 
{21'b111111111111100001000, 21'b000000000000101011001, 21'b000000000000101000101, 21'b111111111111111111110, 21'b111111111111010000011, 21'b111111111111110100100, 21'b111111111111001110111, 21'b111111111111111000111, 21'b000000000000010011000, 21'b111111111111110110011, 21'b111111111111111100000, 21'b111111111111111010111, 21'b111111111111111111111, 21'b111111111111101000100, 21'b111111111111111100100, 21'b111111111111110011001, 21'b000000000000101000000, 21'b111111111111111111111, 21'b111111111110101101111, 21'b000000000000111011100, 21'b000000000001001100001, 21'b000000000000110101000, 21'b111111111111010111011, 21'b111111111111101110011, 21'b111111111111010011101, 21'b111111111111011010111, 21'b000000000000011101000, 21'b000000000000011101111, 21'b000000000000011100111, 21'b000000000000101110000, 21'b000000000000000100011, 21'b000000000000110001011, 21'b111111111111111010101, 21'b000000000000000000100, 21'b000000000000100110111, 21'b000000000000010000110, 21'b111111111111110111100, 21'b111111111111111110110, 21'b000000000000000000000, 21'b111111111111011010100, 21'b111111111111100011011, 21'b111111111111110001111, 21'b111111111111010010000, 21'b000000000000111001100, 21'b000000000000000000000, 21'b111111111111111111010, 21'b111111111111110101011, 21'b111111111111101101000, 21'b111111111110011000111, 21'b111111111111111011000, 21'b111111111111100011010, 21'b111111111111101101110, 21'b111111111111110011001, 21'b000000000000100001110, 21'b000000000001010111010, 21'b000000000000010111111, 21'b111111111111111110010, 21'b111111111111010100000, 21'b111111111111111100001, 21'b000000000000000000000, 21'b000000000000101001101, 21'b111111111111111101010, 21'b000000000000000101110, 21'b000000000000000000000}
};

localparam logic signed [20:0] bias [64] = '{
21'b111111111111111011001,  // -0.037350185215473175
21'b000000000000100011000,  // 0.27355897426605225
21'b111111111111110000001,  // -0.12378914654254913
21'b111111111111110111101,  // -0.064457006752491
21'b000000000000000110111,  // 0.05452875792980194
21'b000000000000001110111,  // 0.11671770364046097
21'b000000000000010001011,  // 0.13640816509723663
21'b000000000000001001100,  // 0.07482525706291199
21'b000000000000000101111,  // 0.04674031585454941
21'b111111111111100110001,  // -0.20146161317825317
21'b111111111111110011010,  // -0.09910125285387039
21'b000000000000010011010,  // 0.15104414522647858
21'b111111111111110010111,  // -0.10221704095602036
21'b111111111111101101010,  // -0.1461549550294876
21'b111111111111110100111,  // -0.08641516417264938
21'b000000000000010101010,  // 0.16613510251045227
21'b111111111111110101010,  // -0.0836295336484909
21'b111111111111111000101,  // -0.05756539851427078
21'b111111111111111011110,  // -0.03229188174009323
21'b111111111111111100010,  // -0.028388574719429016
21'b000000000000010000001,  // 0.1260243058204651
21'b111111111111111011010,  // -0.037064336240291595
21'b000000000000011000110,  // 0.19336333870887756
21'b000000000000000010101,  // 0.02124214917421341
21'b000000000000111111110,  // 0.4985624849796295
21'b000000000000000010000,  // 0.0158411655575037
21'b111111111111110101011,  // -0.08296407759189606
21'b000000000000001110001,  // 0.11056788265705109
21'b000000000000000001100,  // 0.01173810102045536
21'b111111111111110010000,  // -0.10843746364116669
21'b000000000000100011000,  // 0.27439257502555847
21'b000000000000001011110,  // 0.09199801832437515
21'b000000000000100011000,  // 0.27419957518577576
21'b000000000000100010101,  // 0.27063727378845215
21'b111111111111100000001,  // -0.24828937649726868
21'b000000000000001010000,  // 0.07818280160427094
21'b111111111111111111010,  // -0.005749030504375696
21'b000000000000001101111,  // 0.10850494354963303
21'b000000000000010001011,  // 0.13591453433036804
21'b111111111111110000100,  // -0.12088628858327866
21'b111111111111111000101,  // -0.05666546896100044
21'b000000000000001011111,  // 0.09311636537313461
21'b000000000000000111000,  // 0.05477767437696457
21'b000000000000000011110,  // 0.029585206881165504
21'b111111111111011000000,  // -0.31209176778793335
21'b111111111111110101001,  // -0.08465463668107986
21'b111111111111101010100,  // -0.16775836050510406
21'b000000000000010010111,  // 0.14762157201766968
21'b111111111111100001110,  // -0.23618532717227936
21'b000000000000001000010,  // 0.06535740196704865
21'b111111111111101111100,  // -0.12853026390075684
21'b111111111111101110010,  // -0.13802281022071838
21'b111111111111101100100,  // -0.15156887471675873
21'b000000000000001010001,  // 0.07979883998632431
21'b000000000000010111001,  // 0.18141601979732513
21'b111111111111111001000,  // -0.054039113223552704
21'b111111111111111110101,  // -0.010052933357656002
21'b000000000000001000011,  // 0.06611225008964539
21'b000000000000000110011,  // 0.05053366720676422
21'b000000000000000011011,  // 0.026860840618610382
21'b000000000000000100001,  // 0.03283466026186943
21'b000000000000010011111,  // 0.15558314323425293
21'b111111111111011011010,  // -0.2863388657569885
21'b111111111111110100110   // -0.08769102394580841
};
endpackage