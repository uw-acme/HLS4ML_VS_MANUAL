// Width: 11
// NFRAC: 5
package dense_3_11_5;

localparam logic signed [10:0] weights [32][32] = '{ 
{11'b11111111110, 11'b11111110010, 11'b11111110011, 11'b11111111001, 11'b00000001010, 11'b00000000001, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b00000000100, 11'b11111101111, 11'b11111111110, 11'b00000011011, 11'b11111111000, 11'b11111100010, 11'b11111111110, 11'b00000000011, 11'b00000001101, 11'b11111110100, 11'b11111011101, 11'b11111111110, 11'b00000000001, 11'b11111110011, 11'b00000000000, 11'b00000100000, 11'b11111010001, 11'b11111111000, 11'b11111110011, 11'b11111111011, 11'b00000001101, 11'b11111111010}, 
{11'b00000010111, 11'b00000110111, 11'b00000001100, 11'b11111101010, 11'b00000000111, 11'b11111110111, 11'b11111111100, 11'b00000100010, 11'b00000000000, 11'b11111111111, 11'b11111111110, 11'b11111101101, 11'b11111111001, 11'b00000010001, 11'b11110111100, 11'b11111110000, 11'b11111111111, 11'b11111111111, 11'b11111111110, 11'b11111111010, 11'b11111110111, 11'b11111110111, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b11111011101, 11'b00000000000, 11'b00000001111, 11'b11111111101, 11'b11111101001, 11'b00000000000, 11'b00000000001}, 
{11'b11111100000, 11'b00000000101, 11'b00000000000, 11'b00000001010, 11'b11111101011, 11'b00000000000, 11'b00000000000, 11'b11111100101, 11'b00000010001, 11'b11111110111, 11'b11111110111, 11'b11111010000, 11'b11111110110, 11'b00000010000, 11'b00000001000, 11'b11111111111, 11'b11111111100, 11'b11111111111, 11'b11111100101, 11'b00000000000, 11'b00000000011, 11'b00000000010, 11'b00000000110, 11'b00000011100, 11'b00000000001, 11'b11111100110, 11'b00000011000, 11'b00000000000, 11'b00000000101, 11'b11111111111, 11'b00000000000, 11'b00001001000}, 
{11'b00000011010, 11'b11111111111, 11'b11111111001, 11'b00000101001, 11'b00000100111, 11'b00000000000, 11'b00000000010, 11'b00000011010, 11'b11111110011, 11'b11111111111, 11'b11111100101, 11'b00000000011, 11'b00000001000, 11'b11111101000, 11'b00000000010, 11'b11111111010, 11'b11111111111, 11'b11111110100, 11'b00000000001, 11'b00000000001, 11'b00000000000, 11'b11111111101, 11'b00000100110, 11'b00000010101, 11'b00000010101, 11'b00000001111, 11'b00000010101, 11'b00000000000, 11'b11111111100, 11'b00000011100, 11'b00000001111, 11'b11111111010}, 
{11'b00000100000, 11'b11111111101, 11'b11111101001, 11'b11111001111, 11'b00000011110, 11'b00000000000, 11'b11111100101, 11'b11111101101, 11'b11111111101, 11'b11111001100, 11'b11110111001, 11'b00000011110, 11'b00000101010, 11'b00000100001, 11'b11111011011, 11'b11111001110, 11'b00000000000, 11'b11111110110, 11'b00000001100, 11'b00000001000, 11'b11111110011, 11'b11111111111, 11'b00000101110, 11'b11110101000, 11'b00000000101, 11'b11111010101, 11'b00000000100, 11'b11111110000, 11'b11111101100, 11'b11111111111, 11'b00000000100, 11'b00000100101}, 
{11'b00000000010, 11'b11111111101, 11'b11111101100, 11'b11111101111, 11'b00000010111, 11'b00000000000, 11'b11111101110, 11'b11111110111, 11'b11111100100, 11'b11111111011, 11'b11111111111, 11'b00000001010, 11'b00000000000, 11'b00000010110, 11'b11111011111, 11'b11111110111, 11'b00000000101, 11'b11111101101, 11'b11111110011, 11'b11111111111, 11'b00000000000, 11'b00000010011, 11'b00000011101, 11'b11111111111, 11'b11111111111, 11'b00000011001, 11'b11111011100, 11'b11111111111, 11'b11111110000, 11'b11111111101, 11'b11111111111, 11'b00000000000}, 
{11'b00000000100, 11'b11111101010, 11'b00000000110, 11'b11111111101, 11'b11111111111, 11'b00000001001, 11'b11111111001, 11'b11111010100, 11'b11111111111, 11'b11111110010, 11'b11111100010, 11'b00000011110, 11'b00000000000, 11'b00000101011, 11'b00000110101, 11'b00000000000, 11'b11111111111, 11'b11111101011, 11'b11111111100, 11'b00000010001, 11'b11111001111, 11'b00000001001, 11'b00000010100, 11'b00000000001, 11'b00000001001, 11'b00001001111, 11'b11111100110, 11'b11111111010, 11'b11111110011, 11'b00000011111, 11'b11111111100, 11'b11111110101}, 
{11'b11111011001, 11'b00000000001, 11'b11111010111, 11'b00000011011, 11'b00001000001, 11'b00000000111, 11'b00000000000, 11'b00000000011, 11'b11111111111, 11'b00000001000, 11'b00001010011, 11'b11111111111, 11'b00000011000, 11'b00000100111, 11'b00000110001, 11'b00001000011, 11'b00000000000, 11'b11111100001, 11'b00000010101, 11'b11111111111, 11'b11111010111, 11'b11111110001, 11'b00000000000, 11'b11111111010, 11'b11111011111, 11'b00001111000, 11'b11111110001, 11'b00000000000, 11'b00000000000, 11'b00000111000, 11'b00000000101, 11'b00000011001}, 
{11'b00000011011, 11'b11111111110, 11'b00000000000, 11'b11111111101, 11'b00000000101, 11'b11111111101, 11'b11111111111, 11'b00000001010, 11'b00000001101, 11'b11111101110, 11'b00000001000, 11'b00000001011, 11'b00000000000, 11'b00000010101, 11'b11111110001, 11'b11111001100, 11'b00000000000, 11'b11111111111, 11'b11111111110, 11'b11111100000, 11'b11111111111, 11'b00000000000, 11'b11111110011, 11'b11111111111, 11'b11111111001, 11'b00000001001, 11'b00000010111, 11'b11111111000, 11'b11111111100, 11'b11111111101, 11'b00000000001, 11'b11111100110}, 
{11'b11111110100, 11'b00000011000, 11'b00000000000, 11'b00000000000, 11'b00000110010, 11'b00000010100, 11'b11111111111, 11'b11111011100, 11'b00000000111, 11'b11111010011, 11'b11110100110, 11'b11111111111, 11'b00000000000, 11'b00000011011, 11'b00000000111, 11'b00000000000, 11'b11111101010, 11'b00000000000, 11'b00000000000, 11'b00000000011, 11'b00000001111, 11'b11111111110, 11'b11111101000, 11'b00000000000, 11'b11111111111, 11'b00001000101, 11'b00000010100, 11'b11111111111, 11'b11111111011, 11'b00000101010, 11'b11111111101, 11'b11111111010}, 
{11'b11111011110, 11'b00000001011, 11'b11111111101, 11'b11111111111, 11'b11111110000, 11'b11111100111, 11'b00000000011, 11'b00000001001, 11'b11111111111, 11'b11111110101, 11'b11111011011, 11'b00000001100, 11'b00000010011, 11'b00000000000, 11'b00000110101, 11'b11111011100, 11'b00000000110, 11'b11111100110, 11'b00000010010, 11'b11111111111, 11'b11111111101, 11'b00000000100, 11'b00000000111, 11'b00000000000, 11'b11111100000, 11'b00000000001, 11'b11111011100, 11'b11111111101, 11'b11111111111, 11'b00000101011, 11'b11111110011, 11'b00000000000}, 
{11'b11111111111, 11'b00000000111, 11'b00000000000, 11'b00000011001, 11'b11111111000, 11'b11111111101, 11'b00000000011, 11'b11111111111, 11'b11111111101, 11'b00000101001, 11'b00000101100, 11'b00000000000, 11'b11111101010, 11'b11111010011, 11'b11111111100, 11'b00000000000, 11'b00000000000, 11'b11111111011, 11'b11111100001, 11'b00000011000, 11'b00000000000, 11'b00000010111, 11'b11111111111, 11'b00000100011, 11'b00000000111, 11'b00000010011, 11'b00000011101, 11'b11111111100, 11'b11111100110, 11'b11111100011, 11'b11111111111, 11'b11111010101}, 
{11'b11111110001, 11'b11111111111, 11'b00000000111, 11'b11111100101, 11'b00000000101, 11'b11111111111, 11'b11111110010, 11'b11111111111, 11'b11111110111, 11'b00000000010, 11'b00000000100, 11'b11111111011, 11'b00000000001, 11'b00000001100, 11'b11111010111, 11'b11111110000, 11'b00000001110, 11'b11111110100, 11'b00000000000, 11'b11111111110, 11'b00000001100, 11'b00000000000, 11'b11111111110, 11'b00000000010, 11'b00000010001, 11'b11111111001, 11'b00000000000, 11'b11111100011, 11'b11111110011, 11'b11111111111, 11'b00000001011, 11'b00000000000}, 
{11'b11111011110, 11'b00000011010, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b00000001011, 11'b11111111111, 11'b00000110001, 11'b11111111111, 11'b11111111111, 11'b00000001101, 11'b00000000010, 11'b00000000000, 11'b00000000000, 11'b00000000111, 11'b00000010101, 11'b00000001011, 11'b00000001010, 11'b11111111111, 11'b00000010011, 11'b00000000110, 11'b00000000010, 11'b11111111111, 11'b00000010000, 11'b11111111001, 11'b11111101010, 11'b11111111010, 11'b11111111111, 11'b00000000110, 11'b00000000001, 11'b00000001100, 11'b00000011110}, 
{11'b11111111110, 11'b11111100111, 11'b00000000011, 11'b11111111111, 11'b00000111010, 11'b11111110010, 11'b11111011011, 11'b00000000000, 11'b00000000000, 11'b11111111110, 11'b00000000011, 11'b00000011011, 11'b00000010100, 11'b00000000000, 11'b00000000010, 11'b11111110100, 11'b00000000010, 11'b11111111101, 11'b00000000000, 11'b00000000100, 11'b11111111101, 11'b00000000001, 11'b00000010001, 11'b00000000010, 11'b11111111111, 11'b11111100101, 11'b00000001101, 11'b11111111111, 11'b11111111111, 11'b11111111001, 11'b11111111110, 11'b11111111011}, 
{11'b00000000000, 11'b11111111011, 11'b11111110111, 11'b11111110010, 11'b11111011101, 11'b00000100111, 11'b00000000000, 11'b00000001010, 11'b00000010010, 11'b00000000000, 11'b11111111101, 11'b00000011110, 11'b00000001110, 11'b11111101000, 11'b11111110101, 11'b11111111101, 11'b11111100110, 11'b11111111110, 11'b00000000000, 11'b11111111111, 11'b00000001001, 11'b11111110111, 11'b00000000000, 11'b00000000100, 11'b11111111111, 11'b11111101010, 11'b00000001010, 11'b00000000000, 11'b00000000010, 11'b00000000000, 11'b11111101011, 11'b00000000001}, 
{11'b11111110011, 11'b11111110101, 11'b00000000100, 11'b11111111000, 11'b11111111010, 11'b00000000111, 11'b11111111111, 11'b00000000010, 11'b00000001000, 11'b11111111111, 11'b00000000111, 11'b11111110111, 11'b11111111111, 11'b11111111111, 11'b00000000110, 11'b11111111111, 11'b00000011111, 11'b11111111110, 11'b00000001111, 11'b11111110101, 11'b00000001010, 11'b00000000100, 11'b00000000101, 11'b00000000010, 11'b11111111010, 11'b11111101110, 11'b11111101111, 11'b00000000110, 11'b11111111010, 11'b00000000000, 11'b11111111110, 11'b00000001110}, 
{11'b11111111111, 11'b11111100110, 11'b11111100110, 11'b11111111111, 11'b00000101000, 11'b11111111010, 11'b00000000000, 11'b00000011110, 11'b11111110110, 11'b00000000000, 11'b11111100101, 11'b11111100000, 11'b00000011100, 11'b00000001001, 11'b11111111000, 11'b11111101110, 11'b00000001011, 11'b00000000000, 11'b11111110000, 11'b00000000001, 11'b00000000100, 11'b11111111010, 11'b00000010010, 11'b11111000001, 11'b00000000010, 11'b00000001111, 11'b11111111101, 11'b00000000000, 11'b11111110001, 11'b11111111111, 11'b11111110011, 11'b11111111110}, 
{11'b00000001101, 11'b00000010110, 11'b00000100011, 11'b11111110010, 11'b00000011010, 11'b00000010011, 11'b00000000000, 11'b00000011101, 11'b00000010110, 11'b11111111001, 11'b00000101100, 11'b11111101001, 11'b00000100111, 11'b00000011100, 11'b11110111011, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b00000010000, 11'b11111011111, 11'b00000001110, 11'b11111110010, 11'b11111100000, 11'b11111110101, 11'b00000010101, 11'b11111010101, 11'b11111101010, 11'b11111111101, 11'b11111111111, 11'b11111011011, 11'b00000011001, 11'b00000000000}, 
{11'b11111111100, 11'b00000000000, 11'b11111111111, 11'b11111111111, 11'b11111101001, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b11111111110, 11'b11111111101, 11'b00000001000, 11'b11111111111, 11'b00000000101, 11'b11111101010, 11'b00000000110, 11'b11111111111, 11'b00000001001, 11'b00000011100, 11'b11111101001, 11'b00000000011, 11'b11111111001, 11'b00000001000, 11'b00000001100, 11'b11111111010, 11'b11111101111, 11'b00000000001, 11'b00000110101, 11'b11111111110, 11'b11111111111, 11'b00000010100, 11'b00000000000, 11'b00000110111}, 
{11'b11111011110, 11'b00000000010, 11'b11111110010, 11'b00000011000, 11'b00000000111, 11'b11111111101, 11'b11111111111, 11'b11111111111, 11'b11111101100, 11'b11111111101, 11'b00000000000, 11'b11111011100, 11'b00000000000, 11'b11111111101, 11'b11111111111, 11'b11111111111, 11'b11111111000, 11'b00000000000, 11'b00000000000, 11'b00000001010, 11'b00000000001, 11'b00000000000, 11'b00000000000, 11'b11111111111, 11'b00000000000, 11'b00000000001, 11'b00000100101, 11'b11111111111, 11'b11111111111, 11'b11111111101, 11'b00000001011, 11'b11111111110}, 
{11'b11111111111, 11'b11111110110, 11'b00000001101, 11'b00000000010, 11'b11111101000, 11'b00000000000, 11'b00000010010, 11'b11111111111, 11'b00000000000, 11'b11111111001, 11'b00000000111, 11'b00000000001, 11'b00000010100, 11'b11111011100, 11'b11111111001, 11'b11111111110, 11'b00000001101, 11'b11111100111, 11'b00000000001, 11'b11111001111, 11'b11111111110, 11'b11111111000, 11'b11111111101, 11'b00000010010, 11'b11111111011, 11'b11111101110, 11'b00000000101, 11'b00000000000, 11'b00000011001, 11'b00000100001, 11'b11111101011, 11'b11111100011}, 
{11'b00000000100, 11'b00000000001, 11'b11111100101, 11'b11111111100, 11'b11111111111, 11'b00000000000, 11'b00000000110, 11'b00000011010, 11'b00000000000, 11'b00000000001, 11'b00000000100, 11'b11111011101, 11'b11111111011, 11'b11111011001, 11'b00000011110, 11'b00000000000, 11'b11111111111, 11'b11111010110, 11'b11111111111, 11'b11111111011, 11'b11111111110, 11'b00000000000, 11'b00000000011, 11'b11111110110, 11'b00000000011, 11'b00000011010, 11'b00000011011, 11'b00000011000, 11'b00000010011, 11'b00000000000, 11'b00000000111, 11'b00000110010}, 
{11'b11111111110, 11'b11111110000, 11'b00000011000, 11'b11111111001, 11'b00000000100, 11'b00000001010, 11'b11111111111, 11'b11111101101, 11'b11111111010, 11'b11111011001, 11'b00000011100, 11'b00000000000, 11'b00000011010, 11'b00000101010, 11'b11111111000, 11'b11111001000, 11'b11111111001, 11'b00000011110, 11'b11111101101, 11'b11111110010, 11'b00000000011, 11'b00000000000, 11'b11111011101, 11'b11111110011, 11'b11111111101, 11'b11111111000, 11'b00000000111, 11'b00000101101, 11'b00000001111, 11'b11111111111, 11'b00000000101, 11'b00000000001}, 
{11'b00000000010, 11'b00000011101, 11'b00000000000, 11'b00000010010, 11'b00000110101, 11'b11111110101, 11'b11111111111, 11'b11111111101, 11'b00000010010, 11'b11111110011, 11'b11111111111, 11'b00000010101, 11'b00000000000, 11'b00000000001, 11'b11110011110, 11'b11111111010, 11'b00000000000, 11'b00000001100, 11'b11111111111, 11'b00000010011, 11'b11111111111, 11'b11111110100, 11'b11111011100, 11'b00000001000, 11'b00000010010, 11'b11110111001, 11'b11111111111, 11'b00000000000, 11'b00000100010, 11'b11111001100, 11'b00000000000, 11'b11111111111}, 
{11'b00000000000, 11'b11111101010, 11'b00000000011, 11'b11111111111, 11'b00000000011, 11'b00000100001, 11'b11111010001, 11'b00000000010, 11'b00000011011, 11'b11111101010, 11'b11111111110, 11'b00000000011, 11'b11111111111, 11'b00000001011, 11'b00000000110, 11'b11111111110, 11'b00000000100, 11'b00000000000, 11'b00000000001, 11'b00000011000, 11'b11111111110, 11'b11111100001, 11'b11111011001, 11'b11111110011, 11'b11111011010, 11'b00000001101, 11'b00000100111, 11'b00000010111, 11'b11111111111, 11'b11111101000, 11'b11111101100, 11'b00000000011}, 
{11'b00000000011, 11'b11111100001, 11'b11111111110, 11'b00000001001, 11'b11111100001, 11'b00000001010, 11'b11111111111, 11'b11111111111, 11'b11111111111, 11'b00000000000, 11'b00000010000, 11'b11111111110, 11'b00000000000, 11'b00000000000, 11'b00000001000, 11'b11111111110, 11'b00000000000, 11'b11111111111, 11'b11111101011, 11'b11111011111, 11'b11111111111, 11'b11111011101, 11'b11111101100, 11'b11111101000, 11'b00000111000, 11'b00000000001, 11'b11111111101, 11'b00000010100, 11'b00000111001, 11'b00000011001, 11'b11110111100, 11'b11111110100}, 
{11'b00000011000, 11'b11111111111, 11'b00000010000, 11'b11111111110, 11'b00000011110, 11'b11111110110, 11'b00000000100, 11'b00000011010, 11'b00000010001, 11'b11111011110, 11'b11111111100, 11'b00000000111, 11'b00000000100, 11'b11111111111, 11'b00000000101, 11'b00000000000, 11'b00000010111, 11'b00000000010, 11'b00000010111, 11'b11111111011, 11'b11111110111, 11'b11111111011, 11'b11111111111, 11'b00000010011, 11'b11111110011, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b00000000000, 11'b00000010010, 11'b11111101011, 11'b11111111110}, 
{11'b11111111111, 11'b11111111110, 11'b11111100010, 11'b00000010010, 11'b00000001110, 11'b11111111000, 11'b11111111111, 11'b11111110001, 11'b00000000000, 11'b11111111111, 11'b11111101100, 11'b11111110000, 11'b00000011110, 11'b00000000000, 11'b11111110111, 11'b11111111111, 11'b00000001101, 11'b11111111111, 11'b11111111111, 11'b11111110010, 11'b00000010100, 11'b00000000000, 11'b00000001001, 11'b11111111110, 11'b00000001010, 11'b00000000000, 11'b00000000000, 11'b00000001111, 11'b11111110011, 11'b11111111101, 11'b00000001010, 11'b11111111001}, 
{11'b11111111110, 11'b11111101100, 11'b00000100110, 11'b11111111011, 11'b00000001100, 11'b11111101101, 11'b00000000000, 11'b00000000010, 11'b11111100001, 11'b11111111111, 11'b11111111000, 11'b00000000011, 11'b11111101011, 11'b00000001000, 11'b00000001100, 11'b00000000111, 11'b00000000101, 11'b11111111101, 11'b11111010010, 11'b11111111111, 11'b11111111100, 11'b00000001000, 11'b11111111000, 11'b11111111111, 11'b00000001100, 11'b11111111101, 11'b11111111111, 11'b00000011000, 11'b11111100110, 11'b11111101101, 11'b00000010110, 11'b00000000010}, 
{11'b00000011011, 11'b00000001100, 11'b00000000000, 11'b11111110101, 11'b11111111010, 11'b11111111111, 11'b00000000000, 11'b11111111011, 11'b11111111000, 11'b11111111000, 11'b00000000000, 11'b00000001010, 11'b00000000000, 11'b00000000011, 11'b11111111101, 11'b00000000000, 11'b11111110110, 11'b00000000000, 11'b11111111110, 11'b11111111111, 11'b00000000000, 11'b00000000011, 11'b00000000110, 11'b00000000000, 11'b00000000000, 11'b11111011000, 11'b11111110011, 11'b00000000000, 11'b00000000001, 11'b00000000000, 11'b11111110100, 11'b00000000001}, 
{11'b00000001100, 11'b11110111101, 11'b11111111111, 11'b11111111011, 11'b11111110001, 11'b11111111111, 11'b00000000000, 11'b00000100011, 11'b11111111101, 11'b11111111110, 11'b00000000101, 11'b11111010101, 11'b00000000001, 11'b11111100011, 11'b00000101110, 11'b11111111100, 11'b11111110001, 11'b11111011100, 11'b11111111111, 11'b11111010010, 11'b11111001100, 11'b11111111111, 11'b00000000000, 11'b00000000000, 11'b00000001111, 11'b11111111111, 11'b11111101100, 11'b11111111011, 11'b11111111110, 11'b00000000000, 11'b11111111101, 11'b11111010011}
};

localparam logic signed [10:0] bias [32] = '{
11'b00000010000,  // 0.5280959606170654
11'b00000011010,  // 0.8414360880851746
11'b00000001100,  // 0.397830605506897
11'b00000001101,  // 0.4105983078479767
11'b11110001010,  // -3.657735586166382
11'b11111100011,  // -0.8977976441383362
11'b00000110110,  // 1.7051936388015747
11'b11111010111,  // -1.2765135765075684
11'b11111101101,  // -0.5837795734405518
11'b00001010110,  // 2.699671983718872
11'b00000000110,  // 0.2170683741569519
11'b00000011100,  // 0.8814588785171509
11'b11110101011,  // -2.634300947189331
11'b11111000011,  // -1.877297282218933
11'b00000110101,  // 1.6625694036483765
11'b00001010111,  // 2.7459704875946045
11'b11111110000,  // -0.47838035225868225
11'b00000110110,  // 1.6984987258911133
11'b00000011011,  // 0.8548859357833862
11'b00000100000,  // 1.0045719146728516
11'b00000101101,  // 1.4197649955749512
11'b00000011010,  // 0.832463800907135
11'b00000010001,  // 0.5434179306030273
11'b00000011101,  // 0.9277304410934448
11'b11111110101,  // -0.3426123857498169
11'b11111101110,  // -0.5587119460105896
11'b11111101100,  // -0.6208624839782715
11'b11111010111,  // -1.2802538871765137
11'b00000000001,  // 0.05940237268805504
11'b11111100101,  // -0.8213341236114502
11'b00000011100,  // 0.8783953189849854
11'b11111100001   // -0.949700653553009
};
endpackage