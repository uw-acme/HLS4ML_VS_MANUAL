// Width: 17
// NFRAC: 8
package dense_3_17_9;

localparam logic signed [16:0] weights [32][32] = '{ 
{17'b11111111111110011, 17'b11111111110010000, 17'b11111111110011000, 17'b11111111111001111, 17'b00000000001010111, 17'b00000000000001011, 17'b11111111111111100, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000000100000, 17'b11111111101111001, 17'b11111111111110000, 17'b00000000011011000, 17'b11111111111000010, 17'b11111111100010001, 17'b11111111111110110, 17'b00000000000011100, 17'b00000000001101111, 17'b11111111110100110, 17'b11111111011101111, 17'b11111111111110100, 17'b00000000000001100, 17'b11111111110011000, 17'b00000000000000000, 17'b00000000100000011, 17'b11111111010001011, 17'b11111111111000111, 17'b11111111110011100, 17'b11111111111011001, 17'b00000000001101100, 17'b11111111111010111}, 
{17'b00000000010111111, 17'b00000000110111010, 17'b00000000001100110, 17'b11111111101010111, 17'b00000000000111110, 17'b11111111110111010, 17'b11111111111100100, 17'b00000000100010111, 17'b00000000000000001, 17'b11111111111111111, 17'b11111111111110111, 17'b11111111101101001, 17'b11111111111001100, 17'b00000000010001010, 17'b11111110111100100, 17'b11111111110000111, 17'b11111111111111111, 17'b11111111111111101, 17'b11111111111110010, 17'b11111111111010101, 17'b11111111110111101, 17'b11111111110111001, 17'b00000000000000100, 17'b11111111111111111, 17'b11111111111111110, 17'b11111111011101101, 17'b00000000000000011, 17'b00000000001111000, 17'b11111111111101111, 17'b11111111101001111, 17'b00000000000000000, 17'b00000000000001001}, 
{17'b11111111100000011, 17'b00000000000101111, 17'b00000000000000010, 17'b00000000001010010, 17'b11111111101011110, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111100101001, 17'b00000000010001001, 17'b11111111110111100, 17'b11111111110111101, 17'b11111111010000011, 17'b11111111110110000, 17'b00000000010000010, 17'b00000000001000011, 17'b11111111111111111, 17'b11111111111100010, 17'b11111111111111001, 17'b11111111100101111, 17'b00000000000000000, 17'b00000000000011111, 17'b00000000000010001, 17'b00000000000110101, 17'b00000000011100001, 17'b00000000000001001, 17'b11111111100110110, 17'b00000000011000100, 17'b00000000000000000, 17'b00000000000101010, 17'b11111111111111010, 17'b00000000000000000, 17'b00000001001000100}, 
{17'b00000000011010110, 17'b11111111111111111, 17'b11111111111001110, 17'b00000000101001111, 17'b00000000100111010, 17'b00000000000000000, 17'b00000000000010010, 17'b00000000011010000, 17'b11111111110011010, 17'b11111111111111111, 17'b11111111100101101, 17'b00000000000011110, 17'b00000000001000100, 17'b11111111101000000, 17'b00000000000010111, 17'b11111111111010111, 17'b11111111111111111, 17'b11111111110100010, 17'b00000000000001001, 17'b00000000000001110, 17'b00000000000000100, 17'b11111111111101101, 17'b00000000100110001, 17'b00000000010101111, 17'b00000000010101000, 17'b00000000001111111, 17'b00000000010101110, 17'b00000000000000000, 17'b11111111111100001, 17'b00000000011100111, 17'b00000000001111111, 17'b11111111111010011}, 
{17'b00000000100000000, 17'b11111111111101000, 17'b11111111101001110, 17'b11111111001111111, 17'b00000000011110100, 17'b00000000000000000, 17'b11111111100101101, 17'b11111111101101111, 17'b11111111111101000, 17'b11111111001100001, 17'b11111110111001010, 17'b00000000011110010, 17'b00000000101010110, 17'b00000000100001011, 17'b11111111011011001, 17'b11111111001110011, 17'b00000000000000000, 17'b11111111110110111, 17'b00000000001100110, 17'b00000000001000111, 17'b11111111110011111, 17'b11111111111111100, 17'b00000000101110001, 17'b11111110101000000, 17'b00000000000101101, 17'b11111111010101110, 17'b00000000000100001, 17'b11111111110000000, 17'b11111111101100111, 17'b11111111111111111, 17'b00000000000100011, 17'b00000000100101001}, 
{17'b00000000000010110, 17'b11111111111101010, 17'b11111111101100010, 17'b11111111101111010, 17'b00000000010111110, 17'b00000000000000000, 17'b11111111101110000, 17'b11111111110111010, 17'b11111111100100100, 17'b11111111111011111, 17'b11111111111111111, 17'b00000000001010010, 17'b00000000000000000, 17'b00000000010110111, 17'b11111111011111101, 17'b11111111110111110, 17'b00000000000101101, 17'b11111111101101001, 17'b11111111110011010, 17'b11111111111111111, 17'b00000000000000110, 17'b00000000010011001, 17'b00000000011101111, 17'b11111111111111010, 17'b11111111111111111, 17'b00000000011001101, 17'b11111111011100110, 17'b11111111111111111, 17'b11111111110000110, 17'b11111111111101101, 17'b11111111111111110, 17'b00000000000000011}, 
{17'b00000000000100001, 17'b11111111101010101, 17'b00000000000110111, 17'b11111111111101100, 17'b11111111111111100, 17'b00000000001001101, 17'b11111111111001001, 17'b11111111010100101, 17'b11111111111111111, 17'b11111111110010101, 17'b11111111100010110, 17'b00000000011110001, 17'b00000000000000011, 17'b00000000101011110, 17'b00000000110101000, 17'b00000000000000001, 17'b11111111111111111, 17'b11111111101011110, 17'b11111111111100000, 17'b00000000010001011, 17'b11111111001111111, 17'b00000000001001111, 17'b00000000010100111, 17'b00000000000001001, 17'b00000000001001100, 17'b00000001001111100, 17'b11111111100110110, 17'b11111111111010001, 17'b11111111110011110, 17'b00000000011111001, 17'b11111111111100110, 17'b11111111110101001}, 
{17'b11111111011001110, 17'b00000000000001100, 17'b11111111010111101, 17'b00000000011011110, 17'b00000001000001110, 17'b00000000000111011, 17'b00000000000000001, 17'b00000000000011000, 17'b11111111111111111, 17'b00000000001000001, 17'b00000001010011010, 17'b11111111111111111, 17'b00000000011000011, 17'b00000000100111110, 17'b00000000110001001, 17'b00000001000011001, 17'b00000000000000000, 17'b11111111100001011, 17'b00000000010101100, 17'b11111111111111101, 17'b11111111010111001, 17'b11111111110001011, 17'b00000000000000110, 17'b11111111111010101, 17'b11111111011111111, 17'b00000001111000000, 17'b11111111110001111, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000111000100, 17'b00000000000101101, 17'b00000000011001000}, 
{17'b00000000011011000, 17'b11111111111110110, 17'b00000000000000000, 17'b11111111111101001, 17'b00000000000101001, 17'b11111111111101100, 17'b11111111111111111, 17'b00000000001010000, 17'b00000000001101100, 17'b11111111101110011, 17'b00000000001000111, 17'b00000000001011111, 17'b00000000000000110, 17'b00000000010101010, 17'b11111111110001100, 17'b11111111001100111, 17'b00000000000000000, 17'b11111111111111000, 17'b11111111111110010, 17'b11111111100000000, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111110011000, 17'b11111111111111000, 17'b11111111111001111, 17'b00000000001001111, 17'b00000000010111111, 17'b11111111111000010, 17'b11111111111100110, 17'b11111111111101011, 17'b00000000000001101, 17'b11111111100110111}, 
{17'b11111111110100101, 17'b00000000011000100, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000110010101, 17'b00000000010100100, 17'b11111111111111111, 17'b11111111011100011, 17'b00000000000111100, 17'b11111111010011010, 17'b11111110100110001, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000011011011, 17'b00000000000111000, 17'b00000000000000000, 17'b11111111101010111, 17'b00000000000000000, 17'b00000000000000011, 17'b00000000000011111, 17'b00000000001111100, 17'b11111111111110010, 17'b11111111101000111, 17'b00000000000000100, 17'b11111111111111010, 17'b00000001000101001, 17'b00000000010100111, 17'b11111111111111111, 17'b11111111111011011, 17'b00000000101010110, 17'b11111111111101011, 17'b11111111111010011}, 
{17'b11111111011110100, 17'b00000000001011001, 17'b11111111111101110, 17'b11111111111111111, 17'b11111111110000001, 17'b11111111100111110, 17'b00000000000011000, 17'b00000000001001001, 17'b11111111111111111, 17'b11111111110101000, 17'b11111111011011010, 17'b00000000001100110, 17'b00000000010011011, 17'b00000000000000000, 17'b00000000110101101, 17'b11111111011100000, 17'b00000000000110101, 17'b11111111100110111, 17'b00000000010010000, 17'b11111111111111111, 17'b11111111111101100, 17'b00000000000100011, 17'b00000000000111110, 17'b00000000000000000, 17'b11111111100000011, 17'b00000000000001111, 17'b11111111011100001, 17'b11111111111101011, 17'b11111111111111111, 17'b00000000101011001, 17'b11111111110011110, 17'b00000000000000000}, 
{17'b11111111111111111, 17'b00000000000111010, 17'b00000000000000000, 17'b00000000011001000, 17'b11111111111000100, 17'b11111111111101001, 17'b00000000000011101, 17'b11111111111111101, 17'b11111111111101000, 17'b00000000101001000, 17'b00000000101100101, 17'b00000000000000000, 17'b11111111101010101, 17'b11111111010011000, 17'b11111111111100110, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111011111, 17'b11111111100001100, 17'b00000000011000011, 17'b00000000000000001, 17'b00000000010111101, 17'b11111111111111111, 17'b00000000100011111, 17'b00000000000111111, 17'b00000000010011100, 17'b00000000011101001, 17'b11111111111100101, 17'b11111111100110111, 17'b11111111100011110, 17'b11111111111111101, 17'b11111111010101001}, 
{17'b11111111110001100, 17'b11111111111111111, 17'b00000000000111101, 17'b11111111100101001, 17'b00000000000101100, 17'b11111111111111111, 17'b11111111110010000, 17'b11111111111111011, 17'b11111111110111111, 17'b00000000000010011, 17'b00000000000100111, 17'b11111111111011011, 17'b00000000000001000, 17'b00000000001100000, 17'b11111111010111111, 17'b11111111110000010, 17'b00000000001110100, 17'b11111111110100101, 17'b00000000000000000, 17'b11111111111110011, 17'b00000000001100010, 17'b00000000000000100, 17'b11111111111110000, 17'b00000000000010101, 17'b00000000010001001, 17'b11111111111001010, 17'b00000000000000000, 17'b11111111100011000, 17'b11111111110011011, 17'b11111111111111100, 17'b00000000001011000, 17'b00000000000000000}, 
{17'b11111111011110101, 17'b00000000011010111, 17'b11111111111111111, 17'b11111111111111100, 17'b11111111111111011, 17'b00000000001011001, 17'b11111111111111111, 17'b00000000110001011, 17'b11111111111111000, 17'b11111111111111111, 17'b00000000001101001, 17'b00000000000010100, 17'b00000000000000011, 17'b00000000000000000, 17'b00000000000111110, 17'b00000000010101001, 17'b00000000001011011, 17'b00000000001010101, 17'b11111111111111011, 17'b00000000010011101, 17'b00000000000110011, 17'b00000000000010100, 17'b11111111111111011, 17'b00000000010000010, 17'b11111111111001101, 17'b11111111101010010, 17'b11111111111010000, 17'b11111111111111111, 17'b00000000000110100, 17'b00000000000001111, 17'b00000000001100100, 17'b00000000011110101}, 
{17'b11111111111110110, 17'b11111111100111000, 17'b00000000000011010, 17'b11111111111111111, 17'b00000000111010101, 17'b11111111110010101, 17'b11111111011011011, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111110010, 17'b00000000000011000, 17'b00000000011011111, 17'b00000000010100100, 17'b00000000000000101, 17'b00000000000010001, 17'b11111111110100110, 17'b00000000000010001, 17'b11111111111101100, 17'b00000000000000000, 17'b00000000000100110, 17'b11111111111101100, 17'b00000000000001001, 17'b00000000010001000, 17'b00000000000010010, 17'b11111111111111001, 17'b11111111100101100, 17'b00000000001101000, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111001001, 17'b11111111111110101, 17'b11111111111011111}, 
{17'b00000000000000011, 17'b11111111111011111, 17'b11111111110111111, 17'b11111111110010000, 17'b11111111011101000, 17'b00000000100111000, 17'b00000000000000000, 17'b00000000001010110, 17'b00000000010010010, 17'b00000000000000110, 17'b11111111111101110, 17'b00000000011110011, 17'b00000000001110010, 17'b11111111101000100, 17'b11111111110101100, 17'b11111111111101010, 17'b11111111100110100, 17'b11111111111110111, 17'b00000000000000000, 17'b11111111111111101, 17'b00000000001001111, 17'b11111111110111001, 17'b00000000000000000, 17'b00000000000100111, 17'b11111111111111111, 17'b11111111101010001, 17'b00000000001010000, 17'b00000000000000000, 17'b00000000000010110, 17'b00000000000000101, 17'b11111111101011110, 17'b00000000000001010}, 
{17'b11111111110011011, 17'b11111111110101111, 17'b00000000000100111, 17'b11111111111000000, 17'b11111111111010010, 17'b00000000000111011, 17'b11111111111111101, 17'b00000000000010001, 17'b00000000001000011, 17'b11111111111111111, 17'b00000000000111111, 17'b11111111110111110, 17'b11111111111111011, 17'b11111111111111111, 17'b00000000000110100, 17'b11111111111111111, 17'b00000000011111010, 17'b11111111111110111, 17'b00000000001111111, 17'b11111111110101001, 17'b00000000001010001, 17'b00000000000100000, 17'b00000000000101011, 17'b00000000000010010, 17'b11111111111010110, 17'b11111111101110001, 17'b11111111101111011, 17'b00000000000110111, 17'b11111111111010101, 17'b00000000000000000, 17'b11111111111110001, 17'b00000000001110110}, 
{17'b11111111111111111, 17'b11111111100110000, 17'b11111111100110100, 17'b11111111111111111, 17'b00000000101000011, 17'b11111111111010001, 17'b00000000000000000, 17'b00000000011110111, 17'b11111111110110100, 17'b00000000000000000, 17'b11111111100101010, 17'b11111111100000101, 17'b00000000011100101, 17'b00000000001001101, 17'b11111111111000001, 17'b11111111101110011, 17'b00000000001011000, 17'b00000000000000000, 17'b11111111110000110, 17'b00000000000001101, 17'b00000000000100011, 17'b11111111111010010, 17'b00000000010010001, 17'b11111111000001010, 17'b00000000000010100, 17'b00000000001111010, 17'b11111111111101010, 17'b00000000000000111, 17'b11111111110001000, 17'b11111111111111111, 17'b11111111110011001, 17'b11111111111110011}, 
{17'b00000000001101100, 17'b00000000010110000, 17'b00000000100011001, 17'b11111111110010111, 17'b00000000011010101, 17'b00000000010011100, 17'b00000000000000000, 17'b00000000011101001, 17'b00000000010110110, 17'b11111111111001001, 17'b00000000101100111, 17'b11111111101001101, 17'b00000000100111110, 17'b00000000011100100, 17'b11111110111011010, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000000010, 17'b00000000010000101, 17'b11111111011111110, 17'b00000000001110001, 17'b11111111110010011, 17'b11111111100000100, 17'b11111111110101111, 17'b00000000010101000, 17'b11111111010101110, 17'b11111111101010111, 17'b11111111111101010, 17'b11111111111111111, 17'b11111111011011111, 17'b00000000011001010, 17'b00000000000000000}, 
{17'b11111111111100110, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111101001100, 17'b00000000000000100, 17'b00000000000000100, 17'b11111111111111000, 17'b11111111111110011, 17'b11111111111101000, 17'b00000000001000111, 17'b11111111111111111, 17'b00000000000101010, 17'b11111111101010000, 17'b00000000000110110, 17'b11111111111111111, 17'b00000000001001000, 17'b00000000011100101, 17'b11111111101001011, 17'b00000000000011010, 17'b11111111111001101, 17'b00000000001000001, 17'b00000000001100001, 17'b11111111111010100, 17'b11111111101111111, 17'b00000000000001010, 17'b00000000110101000, 17'b11111111111110011, 17'b11111111111111000, 17'b00000000010100110, 17'b00000000000000000, 17'b00000000110111001}, 
{17'b11111111011110100, 17'b00000000000010010, 17'b11111111110010001, 17'b00000000011000100, 17'b00000000000111000, 17'b11111111111101111, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111101100100, 17'b11111111111101111, 17'b00000000000000000, 17'b11111111011100011, 17'b00000000000000110, 17'b11111111111101011, 17'b11111111111111110, 17'b11111111111111111, 17'b11111111111000100, 17'b00000000000000010, 17'b00000000000000001, 17'b00000000001010001, 17'b00000000000001000, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111111111011, 17'b00000000000000000, 17'b00000000000001001, 17'b00000000100101001, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111101011, 17'b00000000001011001, 17'b11111111111110010}, 
{17'b11111111111111111, 17'b11111111110110010, 17'b00000000001101000, 17'b00000000000010100, 17'b11111111101000001, 17'b00000000000000000, 17'b00000000010010010, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111001101, 17'b00000000000111010, 17'b00000000000001001, 17'b00000000010100101, 17'b11111111011100111, 17'b11111111111001111, 17'b11111111111110111, 17'b00000000001101110, 17'b11111111100111011, 17'b00000000000001010, 17'b11111111001111101, 17'b11111111111110110, 17'b11111111111000011, 17'b11111111111101011, 17'b00000000010010111, 17'b11111111111011001, 17'b11111111101110000, 17'b00000000000101110, 17'b00000000000000000, 17'b00000000011001010, 17'b00000000100001011, 17'b11111111101011000, 17'b11111111100011010}, 
{17'b00000000000100010, 17'b00000000000001101, 17'b11111111100101011, 17'b11111111111100010, 17'b11111111111111111, 17'b00000000000000001, 17'b00000000000110110, 17'b00000000011010010, 17'b00000000000000000, 17'b00000000000001010, 17'b00000000000100011, 17'b11111111011101011, 17'b11111111111011101, 17'b11111111011001010, 17'b00000000011110110, 17'b00000000000000000, 17'b11111111111111111, 17'b11111111010110111, 17'b11111111111111111, 17'b11111111111011001, 17'b11111111111110101, 17'b00000000000000000, 17'b00000000000011111, 17'b11111111110110011, 17'b00000000000011011, 17'b00000000011010010, 17'b00000000011011010, 17'b00000000011000111, 17'b00000000010011101, 17'b00000000000000000, 17'b00000000000111010, 17'b00000000110010001}, 
{17'b11111111111110011, 17'b11111111110000110, 17'b00000000011000111, 17'b11111111111001011, 17'b00000000000100011, 17'b00000000001010101, 17'b11111111111111111, 17'b11111111101101101, 17'b11111111111010100, 17'b11111111011001100, 17'b00000000011100101, 17'b00000000000000001, 17'b00000000011010110, 17'b00000000101010111, 17'b11111111111000100, 17'b11111111001000010, 17'b11111111111001010, 17'b00000000011110000, 17'b11111111101101111, 17'b11111111110010101, 17'b00000000000011110, 17'b00000000000000000, 17'b11111111011101000, 17'b11111111110011110, 17'b11111111111101011, 17'b11111111111000001, 17'b00000000000111001, 17'b00000000101101000, 17'b00000000001111101, 17'b11111111111111111, 17'b00000000000101001, 17'b00000000000001110}, 
{17'b00000000000010101, 17'b00000000011101000, 17'b00000000000000000, 17'b00000000010010111, 17'b00000000110101001, 17'b11111111110101000, 17'b11111111111111111, 17'b11111111111101001, 17'b00000000010010110, 17'b11111111110011101, 17'b11111111111111111, 17'b00000000010101010, 17'b00000000000000100, 17'b00000000000001110, 17'b11111110011110010, 17'b11111111111010111, 17'b00000000000000000, 17'b00000000001100110, 17'b11111111111111110, 17'b00000000010011000, 17'b11111111111111111, 17'b11111111110100111, 17'b11111111011100000, 17'b00000000001000010, 17'b00000000010010010, 17'b11111110111001000, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000100010110, 17'b11111111001100101, 17'b00000000000000000, 17'b11111111111111100}, 
{17'b00000000000000100, 17'b11111111101010010, 17'b00000000000011011, 17'b11111111111111000, 17'b00000000000011010, 17'b00000000100001110, 17'b11111111010001100, 17'b00000000000010001, 17'b00000000011011000, 17'b11111111101010011, 17'b11111111111110100, 17'b00000000000011001, 17'b11111111111111011, 17'b00000000001011011, 17'b00000000000110110, 17'b11111111111110111, 17'b00000000000100010, 17'b00000000000000000, 17'b00000000000001011, 17'b00000000011000010, 17'b11111111111110001, 17'b11111111100001000, 17'b11111111011001010, 17'b11111111110011100, 17'b11111111011010001, 17'b00000000001101010, 17'b00000000100111111, 17'b00000000010111100, 17'b11111111111111010, 17'b11111111101000001, 17'b11111111101100000, 17'b00000000000011110}, 
{17'b00000000000011010, 17'b11111111100001011, 17'b11111111111110111, 17'b00000000001001101, 17'b11111111100001011, 17'b00000000001010110, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000010000111, 17'b11111111111110111, 17'b00000000000000100, 17'b00000000000000000, 17'b00000000001000001, 17'b11111111111110111, 17'b00000000000000001, 17'b11111111111111111, 17'b11111111101011011, 17'b11111111011111101, 17'b11111111111111111, 17'b11111111011101110, 17'b11111111101100101, 17'b11111111101000001, 17'b00000000111000111, 17'b00000000000001001, 17'b11111111111101000, 17'b00000000010100010, 17'b00000000111001011, 17'b00000000011001010, 17'b11111110111100001, 17'b11111111110100001}, 
{17'b00000000011000000, 17'b11111111111111111, 17'b00000000010000000, 17'b11111111111110101, 17'b00000000011110111, 17'b11111111110110110, 17'b00000000000100100, 17'b00000000011010110, 17'b00000000010001001, 17'b11111111011110100, 17'b11111111111100000, 17'b00000000000111110, 17'b00000000000100011, 17'b11111111111111000, 17'b00000000000101011, 17'b00000000000000000, 17'b00000000010111001, 17'b00000000000010001, 17'b00000000010111111, 17'b11111111111011110, 17'b11111111110111110, 17'b11111111111011001, 17'b11111111111111111, 17'b00000000010011010, 17'b11111111110011000, 17'b11111111111111100, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000010010101, 17'b11111111101011011, 17'b11111111111110100}, 
{17'b11111111111111111, 17'b11111111111110000, 17'b11111111100010001, 17'b00000000010010001, 17'b00000000001110010, 17'b11111111111000111, 17'b11111111111111111, 17'b11111111110001011, 17'b00000000000000011, 17'b11111111111111111, 17'b11111111101100101, 17'b11111111110000001, 17'b00000000011110101, 17'b00000000000000000, 17'b11111111110111110, 17'b11111111111111111, 17'b00000000001101101, 17'b11111111111111111, 17'b11111111111111111, 17'b11111111110010001, 17'b00000000010100001, 17'b00000000000000000, 17'b00000000001001111, 17'b11111111111110001, 17'b00000000001010000, 17'b00000000000000001, 17'b00000000000000000, 17'b00000000001111011, 17'b11111111110011101, 17'b11111111111101000, 17'b00000000001010010, 17'b11111111111001001}, 
{17'b11111111111110111, 17'b11111111101100010, 17'b00000000100110000, 17'b11111111111011110, 17'b00000000001100100, 17'b11111111101101101, 17'b00000000000000000, 17'b00000000000010001, 17'b11111111100001010, 17'b11111111111111001, 17'b11111111111000000, 17'b00000000000011101, 17'b11111111101011000, 17'b00000000001000110, 17'b00000000001100111, 17'b00000000000111000, 17'b00000000000101011, 17'b11111111111101100, 17'b11111111010010101, 17'b11111111111111001, 17'b11111111111100010, 17'b00000000001000111, 17'b11111111111000111, 17'b11111111111111111, 17'b00000000001100101, 17'b11111111111101000, 17'b11111111111111000, 17'b00000000011000111, 17'b11111111100110100, 17'b11111111101101000, 17'b00000000010110011, 17'b00000000000010010}, 
{17'b00000000011011100, 17'b00000000001100111, 17'b00000000000000000, 17'b11111111110101110, 17'b11111111111010111, 17'b11111111111111111, 17'b00000000000000000, 17'b11111111111011100, 17'b11111111111000000, 17'b11111111111000011, 17'b00000000000000000, 17'b00000000001010001, 17'b00000000000000011, 17'b00000000000011011, 17'b11111111111101001, 17'b00000000000000010, 17'b11111111110110001, 17'b00000000000000000, 17'b11111111111110110, 17'b11111111111111111, 17'b00000000000000001, 17'b00000000000011110, 17'b00000000000110001, 17'b00000000000000000, 17'b00000000000000000, 17'b11111111011000111, 17'b11111111110011001, 17'b00000000000000011, 17'b00000000000001010, 17'b00000000000000000, 17'b11111111110100101, 17'b00000000000001010}, 
{17'b00000000001100000, 17'b11111110111101001, 17'b11111111111111111, 17'b11111111111011001, 17'b11111111110001000, 17'b11111111111111011, 17'b00000000000000000, 17'b00000000100011000, 17'b11111111111101001, 17'b11111111111110100, 17'b00000000000101010, 17'b11111111010101101, 17'b00000000000001100, 17'b11111111100011111, 17'b00000000101110001, 17'b11111111111100101, 17'b11111111110001100, 17'b11111111011100111, 17'b11111111111111010, 17'b11111111010010101, 17'b11111111001100001, 17'b11111111111111111, 17'b00000000000000000, 17'b00000000000000000, 17'b00000000001111100, 17'b11111111111111000, 17'b11111111101100111, 17'b11111111111011010, 17'b11111111111110100, 17'b00000000000000000, 17'b11111111111101111, 17'b11111111010011001}
};

localparam logic signed [16:0] bias [32] = '{
17'b00000000010000111,  // 0.5280959606170654
17'b00000000011010111,  // 0.8414360880851746
17'b00000000001100101,  // 0.397830605506897
17'b00000000001101001,  // 0.4105983078479767
17'b11111110001010111,  // -3.657735586166382
17'b11111111100011010,  // -0.8977976441383362
17'b00000000110110100,  // 1.7051936388015747
17'b11111111010111001,  // -1.2765135765075684
17'b11111111101101010,  // -0.5837795734405518
17'b00000001010110011,  // 2.699671983718872
17'b00000000000110111,  // 0.2170683741569519
17'b00000000011100001,  // 0.8814588785171509
17'b11111110101011101,  // -2.634300947189331
17'b11111111000011111,  // -1.877297282218933
17'b00000000110101001,  // 1.6625694036483765
17'b00000001010111110,  // 2.7459704875946045
17'b11111111110000101,  // -0.47838035225868225
17'b00000000110110010,  // 1.6984987258911133
17'b00000000011011010,  // 0.8548859357833862
17'b00000000100000001,  // 1.0045719146728516
17'b00000000101101011,  // 1.4197649955749512
17'b00000000011010101,  // 0.832463800907135
17'b00000000010001011,  // 0.5434179306030273
17'b00000000011101101,  // 0.9277304410934448
17'b11111111110101000,  // -0.3426123857498169
17'b11111111101110000,  // -0.5587119460105896
17'b11111111101100001,  // -0.6208624839782715
17'b11111111010111000,  // -1.2802538871765137
17'b00000000000001111,  // 0.05940237268805504
17'b11111111100101101,  // -0.8213341236114502
17'b00000000011100000,  // 0.8783953189849854
17'b11111111100001100   // -0.949700653553009
};
endpackage