// Width: 28
// NFRAC: 14
package dense_2_28_14;

localparam logic signed [27:0] weights [64][32] = '{ 
{28'b0000000000000001000100110110, 28'b0000000000000000000010000100, 28'b1111111111111111001111011000, 28'b1111111111111111111010100110, 28'b0000000000000001000010110110, 28'b0000000000000000000000000000, 28'b1111111111111111011011000010, 28'b1111111111111111111111111110, 28'b1111111111111110111001111001, 28'b0000000000000000010100011010, 28'b0000000000000000000000000000, 28'b1111111111111111111110100010, 28'b1111111111111111111111111001, 28'b1111111111111111001100110011, 28'b1111111111111111110011000010, 28'b1111111111111110111100111110, 28'b0000000000000000000000000000, 28'b1111111111111111111100101011, 28'b1111111111111111001111001111, 28'b1111111111111111010111011101, 28'b0000000000000000000000000001, 28'b0000000000000000000000000000, 28'b1111111111111111111101111100, 28'b1111111111111111111111010011, 28'b0000000000000000000000000000, 28'b0000000000000000011001101110, 28'b0000000000000001100010110101, 28'b0000000000000000101100110111, 28'b1111111111111111111111111000, 28'b0000000000000000001100111101, 28'b1111111111111110010111001101, 28'b0000000000000000000000000101}, 
{28'b1111111111111111100110010110, 28'b1111111111111111011000010110, 28'b1111111111111111011100100101, 28'b1111111111111111110001110011, 28'b1111111111111111111110100011, 28'b0000000000000000001011000000, 28'b1111111111111111000110110101, 28'b0000000000000000000001010110, 28'b0000000000000000000001001110, 28'b1111111111111111101111111001, 28'b0000000000000000100111111110, 28'b1111111111111111110100111001, 28'b1111111111111111110000111011, 28'b1111111111111111001000011110, 28'b0000000000000000000001111010, 28'b1111111111111111110011101101, 28'b0000000000000000000011001100, 28'b1111111111111111001110001001, 28'b0000000000000000101011111110, 28'b0000000000000000111010110001, 28'b1111111111111111110111111110, 28'b1111111111111111111110100011, 28'b1111111111111111111111111011, 28'b0000000000000000000110000011, 28'b1111111111111111101101110000, 28'b0000000000000001000110011010, 28'b0000000000000000111111011000, 28'b0000000000000000000010001011, 28'b0000000000000000000111010011, 28'b1111111111111110000011011001, 28'b0000000000000000000001111000, 28'b0000000000000000000000000000}, 
{28'b0000000000000000010010100011, 28'b1111111111111111100010101000, 28'b1111111111111111011110110100, 28'b1111111111111111110101010011, 28'b1111111111111111101100001011, 28'b1111111111111111101010001010, 28'b1111111111111111010000101010, 28'b0000000000000000000001001001, 28'b1111111111111111011101011100, 28'b0000000000000000000010010010, 28'b0000000000000000000000100010, 28'b1111111111111111101011010110, 28'b0000000000000000010111001001, 28'b1111111111111111101111011111, 28'b1111111111111111111111101001, 28'b1111111111111111110110100110, 28'b0000000000000000000001010000, 28'b0000000000000000011000011100, 28'b0000000000000000001111000000, 28'b0000000000000000111010110101, 28'b0000000000000000001010100001, 28'b1111111111111111101010011110, 28'b0000000000000000000000000110, 28'b0000000000000000001000111100, 28'b1111111111111111111011010011, 28'b0000000000000000110101100101, 28'b0000000000000000100110001100, 28'b0000000000000000011000110011, 28'b1111111111111111111111111001, 28'b1111111111111111011001000100, 28'b1111111111111111111100100010, 28'b0000000000000000011001011011}, 
{28'b0000000000000000100011010111, 28'b0000000000000000000100111010, 28'b0000000000000000001101100011, 28'b1111111111111111111101100001, 28'b1111111111111101111101101011, 28'b0000000000000000000000000000, 28'b0000000000000000000000000101, 28'b0000000000000000111001111001, 28'b0000000000000000111110000110, 28'b1111111111111111111100100110, 28'b1111111111111111111111111111, 28'b0000000000000000000000000001, 28'b0000000000000000000000000101, 28'b0000000000000000000001010000, 28'b1111111111111111111011010100, 28'b0000000000000000110110111110, 28'b0000000000000000000000000010, 28'b1111111111111111111001101101, 28'b1111111111111111111111111111, 28'b1111111111111111010010111010, 28'b1111111111111111110000010101, 28'b0000000000000000001100101011, 28'b1111111111111111101111110000, 28'b1111111111111111111111111010, 28'b0000000000000000000000111111, 28'b1111111111111111110011000000, 28'b0000000000000000010010101100, 28'b1111111111111111111111111101, 28'b1111111111111111111111111110, 28'b1111111111111111111111111111, 28'b1111111111111111001000111011, 28'b0000000000000001001111011011}, 
{28'b1111111111111101010001010011, 28'b1111111111111111111001101001, 28'b1111111111111111111110111011, 28'b0000000000000000000001010110, 28'b1111111111111111111001010001, 28'b0000000000000000000001101100, 28'b1111111111111111110011011011, 28'b1111111111111111011001101011, 28'b0000000000000000001101111000, 28'b1111111111111111111010110101, 28'b1111111111111111111100100000, 28'b1111111111111111111111111101, 28'b1111111111111111111111111101, 28'b0000000000000000110101110100, 28'b0000000000000000000000000001, 28'b0000000000000001010100001111, 28'b1111111111111111111111111110, 28'b0000000000000000110111110111, 28'b1111111111111110011001100110, 28'b0000000000000000000000000100, 28'b1111111111111111100011011011, 28'b0000000000000000101011001001, 28'b0000000000000001000010000110, 28'b0000000000000000000000000001, 28'b0000000000000000001011100110, 28'b0000000000000000101001101101, 28'b0000000000000000111101000111, 28'b0000000000000000000100011100, 28'b1111111111111111111110110110, 28'b1111111111111111111111111101, 28'b1111111111111111111100011110, 28'b0000000000000000111001111010}, 
{28'b0000000000000000001110110001, 28'b1111111111111111111111111101, 28'b0000000000000000100110001101, 28'b1111111111111101011001111111, 28'b1111111111111010011111011100, 28'b1111111111111110100110010010, 28'b0000000000000001011010101011, 28'b1111111111111101100000101111, 28'b1111111111111111111111111010, 28'b1111111111111101010010100110, 28'b1111111111111101111111101111, 28'b1111111111111110101000101100, 28'b0000000000000001011010011101, 28'b1111111111111111111111111111, 28'b1111111111111111111100001100, 28'b0000000000000000000000000000, 28'b1111111111111111111111111111, 28'b1111111111111111111111111001, 28'b1111111111111111011110001001, 28'b1111111111111111111111111110, 28'b1111111111111110000010110000, 28'b0000000000000000000000000000, 28'b0000000000000000101111100110, 28'b1111111111111111111111111110, 28'b0000000000000000000101101000, 28'b0000000000000001000100100010, 28'b0000000000000000001101000111, 28'b1111111111111111111111111111, 28'b1111111111111111111111111110, 28'b0000000000000000110100101000, 28'b1111111111111111110111010000, 28'b0000000000000000110011010110}, 
{28'b1111111111111111110110110010, 28'b1111111111111111010111101111, 28'b1111111111111111000010001001, 28'b1111111111111111110011111110, 28'b1111111111111110110110001000, 28'b0000000000000000010000111011, 28'b1111111111111111010001111011, 28'b1111111111111111011011101001, 28'b1111111111111110010101110100, 28'b0000000000000000001100011001, 28'b1111111111111111111110101100, 28'b1111111111111111010111010000, 28'b0000000000000000011110011101, 28'b1111111111111111111101011010, 28'b1111111111111111110101011000, 28'b1111111111111101110010010000, 28'b1111111111111111111111111100, 28'b0000000000000000010101100000, 28'b0000000000000000110001000100, 28'b1111111111111111010110011101, 28'b1111111111111111011001100111, 28'b1111111111111111101111111110, 28'b1111111111111111111111101010, 28'b0000000000000000000111000100, 28'b1111111111111111110100010111, 28'b1111111111111101011010000100, 28'b1111111111111110111100001011, 28'b1111111111111111110100011111, 28'b0000000000000000000001011101, 28'b1111111111111111111010100011, 28'b0000000000000000000111110101, 28'b1111111111111111111111110100}, 
{28'b1111111111111111011000101100, 28'b1111111111111111101000110110, 28'b1111111111111111101011101010, 28'b1111111111111111000011010001, 28'b1111111111111111100010010110, 28'b1111111111111111111111111011, 28'b0000000000000000011010101111, 28'b1111111111111111101011110000, 28'b0000000000000000110011010110, 28'b0000000000000000000000000010, 28'b0000000000000000000000000001, 28'b1111111111111111111111111110, 28'b0000000000000000111000000001, 28'b0000000000000000000000000010, 28'b1111111111111111111111111100, 28'b1111111111111111101101111000, 28'b1111111111111111111111111001, 28'b0000000000000000000000000000, 28'b1111111111111111111111111001, 28'b0000000000000000000000000001, 28'b1111111111111111111111111010, 28'b1111111111111111111111110111, 28'b0000000000000000000000000011, 28'b1111111111111111111111111111, 28'b0000000000000000001011010011, 28'b1111111111111111010001111011, 28'b0000000000000000000011100011, 28'b1111111111111111111111111011, 28'b1111111111111111101101100010, 28'b1111111111111111111111110100, 28'b0000000000000000000000000111, 28'b1111111111111111111111111101}, 
{28'b1111111111111110000101110001, 28'b1111111111111111110001011000, 28'b1111111111111110011110101100, 28'b0000000000000000011111010011, 28'b0000000000000001111100101010, 28'b1111111111111111111111111111, 28'b1111111111111111111000100100, 28'b0000000000000000111101001010, 28'b1111111111111110001111101011, 28'b1111111111111111110100000010, 28'b0000000000000000000000000001, 28'b1111111111111111001100011011, 28'b1111111111111111111111111010, 28'b0000000000000000010011011111, 28'b1111111111111111001111001110, 28'b0000000000000011000001000000, 28'b1111111111111111111101110011, 28'b0000000000000000001011111110, 28'b0000000000000000110101001011, 28'b0000000000000000111110101100, 28'b0000000000000000000000000011, 28'b1111111111111110101010000010, 28'b0000000000000000000000000011, 28'b0000000000000001101001010111, 28'b1111111111111111010001100111, 28'b0000000000000010110010100110, 28'b1111111111111111011001110010, 28'b1111111111111111001011110011, 28'b1111111111111110000111001011, 28'b1111111111111110001001001011, 28'b0000000000000000000000000100, 28'b0000000000000000001101101011}, 
{28'b0000000000000000000000000010, 28'b1111111111111111111100000010, 28'b1111111111111111101101000110, 28'b0000000000000000000000000000, 28'b0000000000000001001110111110, 28'b1111111111111111111010110101, 28'b1111111111111111101111101101, 28'b0000000000000000010111100000, 28'b0000000000000000011001111110, 28'b0000000000000000000000111000, 28'b1111111111111111111101110100, 28'b1111111111111111111111111010, 28'b1111111111111111111111111111, 28'b1111111111111111100010111010, 28'b1111111111111111111111111110, 28'b0000000000000000000000000100, 28'b0000000000000000000000000000, 28'b1111111111111111111110101101, 28'b0000000000000000000000100011, 28'b0000000000000000010101101111, 28'b0000000000000000000100111011, 28'b1111111111111111111111111110, 28'b0000000000000000000000000011, 28'b0000000000000000000001110101, 28'b0000000000000000001001110100, 28'b1111111111111111011110001100, 28'b0000000000000000010001011001, 28'b0000000000000000111111101000, 28'b1111111111111111111111111111, 28'b0000000000000000000001100100, 28'b0000000000000000001100101100, 28'b0000000000000000010001110001}, 
{28'b0000000000000000011000101001, 28'b0000000000000000000000000000, 28'b1111111111111111100101100111, 28'b1111111111111110111111110010, 28'b1111111111111100110100101110, 28'b0000000000000000100010000100, 28'b0000000000000000000000000111, 28'b1111111111111100101100001100, 28'b0000000000000000001001010011, 28'b1111111111111111111111111011, 28'b0000000000000000000000111100, 28'b1111111111111111111111100101, 28'b0000000000000000000010101101, 28'b0000000000000000000000000011, 28'b1111111111111111111011001010, 28'b1111111111111110011110010010, 28'b1111111111111111111111111110, 28'b0000000000000000111000010010, 28'b0000000000000000100000010110, 28'b0000000000000000110000111101, 28'b1111111111111110001111011101, 28'b1111111111111110100100111001, 28'b0000000000000000011110101111, 28'b1111111111111111110111000101, 28'b1111111111111111110100001100, 28'b0000000000000001011011110010, 28'b1111111111111111100111010000, 28'b1111111111111111111111111011, 28'b1111111111111111111111111101, 28'b0000000000000000110110000010, 28'b1111111111111111111111111101, 28'b0000000000000000000001100111}, 
{28'b1111111111111111001101011111, 28'b1111111111111110000001110010, 28'b0000000000000000000000000000, 28'b1111111111111111111111011101, 28'b0000000000000001010101000000, 28'b1111111111111110111011000101, 28'b1111111111111111000111010100, 28'b0000000000000000011101101011, 28'b1111111111111111111111110110, 28'b0000000000000000100110000101, 28'b0000000000000000010010111100, 28'b1111111111111111101100101000, 28'b0000000000000000000000000100, 28'b0000000000000000000011100111, 28'b1111111111111111111010100100, 28'b1111111111111110111111001110, 28'b0000000000000000101100111010, 28'b0000000000000000000111010011, 28'b0000000000000001001100000110, 28'b0000000000000000010110001001, 28'b0000000000000000000000000000, 28'b1111111111111111110110010100, 28'b0000000000000000100000010001, 28'b1111111111111111101001111000, 28'b1111111111111110110001001001, 28'b1111111111111111111110010010, 28'b0000000000000000101111010111, 28'b1111111111111111111111111100, 28'b0000000000000000000010001010, 28'b1111111111111111100111110000, 28'b0000000000000000100011001100, 28'b0000000000000001000110101110}, 
{28'b0000000000000000000011111000, 28'b0000000000000000000000000010, 28'b0000000000000000111000001000, 28'b0000000000000000000010001001, 28'b1111111111111111110101100101, 28'b0000000000000000101110001100, 28'b0000000000000000010111100111, 28'b1111111111111111111111111011, 28'b0000000000000000000000001101, 28'b1111111111111111011100000111, 28'b1111111111111111110010000000, 28'b1111111111111111010101001010, 28'b1111111111111111111111111100, 28'b0000000000000000001100111010, 28'b1111111111111111101110010110, 28'b0000000000000011010111110110, 28'b0000000000000000000000000100, 28'b1111111111111111100111111010, 28'b1111111111111111001111101100, 28'b1111111111111111111100100111, 28'b0000000000000000110010110111, 28'b0000000000000000100000110000, 28'b0000000000000000000000000011, 28'b1111111111111111111111010110, 28'b0000000000000000111000001100, 28'b0000000000000001000100101001, 28'b0000000000000001111110110011, 28'b0000000000000000000010101001, 28'b0000000000000000000000000010, 28'b0000000000000000000000000111, 28'b1111111111111111111100111100, 28'b1111111111111111101101101100}, 
{28'b1111111111111111011000000001, 28'b0000000000000000001100011000, 28'b0000000000000000001010000101, 28'b1111111111111111000000101101, 28'b1111111111111110111011000000, 28'b0000000000000001111000000011, 28'b0000000000000000001100100101, 28'b0000000000000000000000000000, 28'b1111111111111111010110110110, 28'b1111111111111111101001011001, 28'b0000000000000000100001001010, 28'b0000000000000000010010001000, 28'b0000000000000000000000001001, 28'b1111111111111111101011111010, 28'b0000000000000001001001001111, 28'b1111111111111111111111111100, 28'b1111111111111111111100100001, 28'b0000000000000000000000000010, 28'b0000000000000000000011010111, 28'b1111111111111111110100000110, 28'b0000000000000000010100000010, 28'b0000000000000000000100000010, 28'b0000000000000000011101001101, 28'b1111111111111111111111111011, 28'b0000000000000000000000110110, 28'b0000000000000010101000011110, 28'b1111111111111111110001100100, 28'b1111111111111111111010000111, 28'b1111111111111111111111111101, 28'b1111111111111111100100000010, 28'b1111111111111111110101101111, 28'b0000000000000000101101000010}, 
{28'b0000000000000000001111000101, 28'b0000000000000000010010111111, 28'b0000000000000001010011100101, 28'b1111111111111111110101110100, 28'b0000000000000000011001110110, 28'b0000000000000001011001110100, 28'b0000000000000000000000001011, 28'b1111111111111111111000011110, 28'b0000000000000000011110001101, 28'b1111111111111111100010110110, 28'b1111111111111111111111111110, 28'b1111111111111111100001011111, 28'b0000000000000000000000000101, 28'b0000000000000001100100101010, 28'b1111111111111111111011011110, 28'b0000000000000000000000011010, 28'b0000000000000000111100011101, 28'b0000000000000000000000001010, 28'b0000000000000000000000110000, 28'b1111111111111110101111111010, 28'b1111111111111111000001001001, 28'b1111111111111111110110110000, 28'b1111111111111111111111111111, 28'b1111111111111111011010101001, 28'b1111111111111111110110110000, 28'b1111111111111111101010111001, 28'b1111111111111111001101101110, 28'b1111111111111111001001100111, 28'b0000000000000000000111101100, 28'b0000000000000000011100100100, 28'b1111111111111110011010010011, 28'b0000000000000000000000110101}, 
{28'b1111111111111110110011100101, 28'b0000000000000000000000000001, 28'b1111111111111111111100001100, 28'b1111111111111111110011010010, 28'b1111111111111111111111111100, 28'b0000000000000000100010001000, 28'b1111111111111111101100001100, 28'b0000000000000001000101011000, 28'b1111111111111110100011000010, 28'b1111111111111111111111110110, 28'b0000000000000000000000000000, 28'b1111111111111111111111111111, 28'b0000000000000000000000000101, 28'b0000000000000000000000000010, 28'b1111111111111111111111000011, 28'b1111111111111111101000110011, 28'b0000000000000000010100010010, 28'b0000000000000000101110111010, 28'b1111111111111111111101100111, 28'b1111111111111110111111101011, 28'b1111111111111111110000111101, 28'b0000000000000000011100101000, 28'b0000000000000000010000001000, 28'b0000000000000000000000000111, 28'b0000000000000000000000110001, 28'b0000000000000000010100111010, 28'b1111111111111111000010101100, 28'b0000000000000000000000000001, 28'b1111111111111111111111111111, 28'b0000000000000000000000110110, 28'b0000000000000000000000001000, 28'b1111111111111111011111110011}, 
{28'b1111111111111110101001111100, 28'b1111111111111111111110100000, 28'b1111111111111111111111001111, 28'b1111111111111111111011100011, 28'b1111111111111111111110110001, 28'b0000000000000000011011000000, 28'b0000000000000000000001101100, 28'b0000000000000000001000110111, 28'b0000000000000000001001110001, 28'b0000000000000000010000000111, 28'b0000000000000000010100001100, 28'b0000000000000000101001010000, 28'b0000000000000000000110110111, 28'b1111111111111111100111001111, 28'b0000000000000000000000001000, 28'b0000000000000001100001101001, 28'b0000000000000000000000000101, 28'b0000000000000000000000010010, 28'b1111111111111111111111010110, 28'b0000000000000000011100001010, 28'b0000000000000000100100011100, 28'b0000000000000000000111111001, 28'b0000000000000000001010100011, 28'b1111111111111111111000011001, 28'b1111111111111111110111110000, 28'b0000000000000000000110110010, 28'b1111111111111111101110110101, 28'b1111111111111111011111100100, 28'b0000000000000000110101101000, 28'b1111111111111111111000001000, 28'b0000000000000000001000000110, 28'b1111111111111111001111111011}, 
{28'b0000000000000000000000000010, 28'b1111111111111111111111111111, 28'b0000000000000000001001101001, 28'b0000000000000000000000000010, 28'b0000000000000011101000000111, 28'b1111111111111111111111110011, 28'b0000000000000000000000000000, 28'b1111111111111111111111111111, 28'b0000000000000000011100000100, 28'b1111111111111111101100110001, 28'b0000000000000000000000000000, 28'b0000000000000000000000000001, 28'b0000000000000000000000010010, 28'b0000000000000000100001000011, 28'b0000000000000000000000000000, 28'b1111111111111111011010110010, 28'b1111111111111111111111111110, 28'b1111111111111111101110110110, 28'b0000000000000001010011110100, 28'b0000000000000000000000000011, 28'b1111111111111111111111111111, 28'b1111111111111111111111111011, 28'b0000000000000000000000000001, 28'b1111111111111111111111111111, 28'b0000000000000000000000000000, 28'b0000000000000000010001011111, 28'b0000000000000000000000000000, 28'b0000000000000000000000000000, 28'b1111111111111111111111111111, 28'b1111111111111111111111111101, 28'b0000000000000000000000000011, 28'b0000000000000000001010100110}, 
{28'b1111111111111111111111001001, 28'b0000000000000000000111011011, 28'b1111111111111111111111110011, 28'b0000000000000000001100010000, 28'b1111111111111111110100101000, 28'b1111111111111111100001011101, 28'b1111111111111111110000000001, 28'b0000000000000001000111000111, 28'b0000000000000000000000000100, 28'b0000000000000000011000110011, 28'b1111111111111111111101001011, 28'b0000000000000000010000100111, 28'b1111111111111111110111100000, 28'b1111111111111111010111101010, 28'b1111111111111111001111001110, 28'b0000000000000000000011010110, 28'b1111111111111111111111111111, 28'b1111111111111111110111000101, 28'b0000000000000000000000000001, 28'b0000000000000000000000000110, 28'b1111111111111111111111110111, 28'b0000000000000000010011011000, 28'b0000000000000000001001001000, 28'b1111111111111111011111110011, 28'b0000000000000000011100100111, 28'b1111111111111111010101111001, 28'b0000000000000000000000100011, 28'b0000000000000000000000000000, 28'b1111111111111111010101000101, 28'b0000000000000000000000000000, 28'b0000000000000000001011101011, 28'b1111111111111111111000000010}, 
{28'b1111111111111111111101000011, 28'b1111111111111111100110101010, 28'b0000000000000000000000000011, 28'b1111111111111111110000101100, 28'b0000000000000000110111010010, 28'b1111111111111111111111111011, 28'b1111111111111111111010101010, 28'b0000000000000000011011010101, 28'b1111111111111110011011111100, 28'b0000000000000000000000000010, 28'b1111111111111111110110001000, 28'b1111111111111111111111011101, 28'b0000000000000001011001111111, 28'b0000000000000000111010101111, 28'b1111111111111111100110100101, 28'b1111111111111111111010101011, 28'b1111111111111111111111111011, 28'b0000000000000000000000001011, 28'b1111111111111111111111111101, 28'b0000000000000000000000000101, 28'b0000000000000000000000000011, 28'b1111111111111111011101001111, 28'b1111111111111111100001100011, 28'b0000000000000000100001100000, 28'b0000000000000000000000000000, 28'b1111111111111111011100111010, 28'b0000000000000000000110010000, 28'b1111111111111111101011011011, 28'b1111111111111111110111011110, 28'b0000000000000000100010110011, 28'b0000000000000000000000001001, 28'b1111111111111111000000101111}, 
{28'b0000000000000010100010011111, 28'b0000000000000001010111100010, 28'b1111111111111111000000001011, 28'b0000000000000000000000110101, 28'b1111111111111110100111011010, 28'b0000000000000000000000000001, 28'b0000000000000000111001000010, 28'b0000000000000000000111111101, 28'b0000000000000000111001010010, 28'b1111111111111111111111111011, 28'b1111111111111111011000010111, 28'b1111111111111111101011111001, 28'b0000000000000000100100010010, 28'b0000000000000000000111000101, 28'b1111111111111111100110110111, 28'b0000000000000000100001101110, 28'b0000000000000010001001000001, 28'b1111111111111111011110101101, 28'b1111111111111110110100001100, 28'b0000000000000000000000000001, 28'b1111111111111111111000101010, 28'b1111111111111111010010110010, 28'b1111111111111111111100111001, 28'b1111111111111111111111100111, 28'b0000000000000000010110000000, 28'b1111111111111110100011101111, 28'b0000000000000000010110110000, 28'b1111111111111111111111101110, 28'b0000000000000000000000000101, 28'b0000000000000000011011111010, 28'b1111111111111111111000100111, 28'b0000000000000000001111010000}, 
{28'b1111111111111111101000010011, 28'b1111111111111111001110110111, 28'b1111111111111111110110101101, 28'b1111111111111111010101001010, 28'b1111111111111111111011100110, 28'b0000000000000000001100100110, 28'b0000000000000000000000000011, 28'b1111111111111111111101000110, 28'b0000000000000000001001101000, 28'b1111111111111111111111000111, 28'b0000000000000000000000000011, 28'b1111111111111111001000011101, 28'b0000000000000000011010000111, 28'b0000000000000000010100100100, 28'b1111111111111111100101110011, 28'b0000000000000001110001100010, 28'b1111111111111111111111111100, 28'b0000000000000000000000000011, 28'b1111111111111111111110111110, 28'b0000000000000000000000000001, 28'b0000000000000001010000111010, 28'b1111111111111110000111100001, 28'b1111111111111111100100010001, 28'b1111111111111111110001101011, 28'b1111111111111111111011001111, 28'b0000000000000000110010011101, 28'b1111111111111111110010100101, 28'b0000000000000000000100100000, 28'b0000000000000001111011111110, 28'b1111111111111101111100110011, 28'b1111111111111110100010000000, 28'b0000000000000000000101101111}, 
{28'b0000000000000000000100010011, 28'b1111111111111111110000111100, 28'b1111111111111111111111111111, 28'b0000000000000000000000000011, 28'b1111111111111101000111111101, 28'b1111111111111101100100110000, 28'b0000000000000000000000011000, 28'b1111111111111111111111111101, 28'b1111111111111110111100001001, 28'b0000000000000000000110010100, 28'b0000000000000000000000000000, 28'b1111111111111111111000111101, 28'b0000000000000000000000000000, 28'b1111111111111111110001000011, 28'b1111111111111111110010100010, 28'b1111111111111111101110010111, 28'b1111111111111111011010010111, 28'b0000000000000001001000010000, 28'b0000000000000000000000000001, 28'b0000000000000000001011110100, 28'b1111111111111111111111111000, 28'b1111111111111111101101111100, 28'b0000000000000000000000000001, 28'b1111111111111111101001110010, 28'b0000000000000000111000001101, 28'b1111111111111101100000101010, 28'b0000000000000000111000010110, 28'b1111111111111111111111111110, 28'b1111111111111111111110110000, 28'b0000000000000000110011001101, 28'b1111111111111111111111111110, 28'b0000000000000000111100011111}, 
{28'b1111111111111111111111111101, 28'b0000000000000000000001010100, 28'b1111111111111111110100111101, 28'b0000000000000000010011001111, 28'b0000000000000000001110001010, 28'b1111111111111110101000011101, 28'b0000000000000000000000000011, 28'b0000000000000000010000011111, 28'b0000000000000010010100011000, 28'b1111111111111111111101101101, 28'b0000000000000000000000000000, 28'b0000000000000000001110011011, 28'b0000000000000001011011111001, 28'b1111111111111111110111110111, 28'b0000000000000000000011100101, 28'b0000000000000000011001110111, 28'b1111111111111111111111111110, 28'b0000000000000000000111000111, 28'b1111111111111111111111111011, 28'b0000000000000000000000001111, 28'b1111111111111110111001111011, 28'b0000000000000000001001110100, 28'b0000000000000000010001111111, 28'b0000000000000000000101110100, 28'b1111111111111111111111111101, 28'b0000000000000000110111111000, 28'b0000000000000000000001001001, 28'b0000000000000000100000010001, 28'b1111111111111110010101000110, 28'b0000000000000000011010010100, 28'b0000000000000001100101010010, 28'b0000000000000000000001011100}, 
{28'b1111111111111110100110001010, 28'b0000000000000000110110000010, 28'b1111111111111110111101010101, 28'b0000000000000000011111011110, 28'b1111111111111111100101000000, 28'b0000000000000000000000000100, 28'b0000000000000001111111011001, 28'b1111111111111111000100011010, 28'b1111111111111110110101011101, 28'b0000000000000000101011110111, 28'b1111111111111111000110111111, 28'b1111111111111111111001111110, 28'b1111111111111111111111110001, 28'b0000000000000001011000000100, 28'b1111111111111111111111100110, 28'b1111111111111110110010110000, 28'b1111111111111111111111111110, 28'b0000000000000001110000110111, 28'b1111111111111110000111011011, 28'b1111111111111111111001110010, 28'b0000000000000001010001000011, 28'b1111111111111110100011001010, 28'b0000000000000000001101100100, 28'b1111111111111111111100001000, 28'b0000000000000001000101011111, 28'b1111111111111101111101110010, 28'b1111111111111110100011001000, 28'b1111111111111111001101110010, 28'b1111111111111111111111111110, 28'b0000000000000000011010100000, 28'b0000000000000000000110011011, 28'b0000000000000000101101101010}, 
{28'b1111111111111111101000110001, 28'b0000000000000000001101010011, 28'b1111111111111111111111111101, 28'b0000000000000000100110010110, 28'b1111111111111111110110010010, 28'b0000000000000000111010000111, 28'b0000000000000000000000100000, 28'b1111111111111111111101001000, 28'b1111111111111111111111011110, 28'b0000000000000000000000010010, 28'b0000000000000000000000000001, 28'b1111111111111111111111111111, 28'b1111111111111111111111100001, 28'b0000000000000010000101001010, 28'b0000000000000000000011001110, 28'b0000000000000000110000010110, 28'b0000000000000000000000000100, 28'b1111111111111111001001110100, 28'b1111111111111111101100011101, 28'b1111111111111111111111111110, 28'b1111111111111111111011110000, 28'b0000000000000000001010110010, 28'b1111111111111111111111111110, 28'b1111111111111111010000100101, 28'b1111111111111111111111111110, 28'b0000000000000001001011101011, 28'b0000000000000001001111011011, 28'b1111111111111111111111111111, 28'b1111111111111111111011110100, 28'b0000000000000000000000000000, 28'b1111111111111111111111110111, 28'b1111111111111111100111010100}, 
{28'b1111111111111111101011010100, 28'b0000000000000000000000000001, 28'b0000000000000001000101111000, 28'b0000000000000000000000000001, 28'b0000000000000000000000000001, 28'b1111111111111111100010111011, 28'b0000000000000000000000000101, 28'b1111111111111100100010111000, 28'b0000000000000000110111001011, 28'b0000000000000000000011100001, 28'b0000000000000000000110110101, 28'b1111111111111110100011111000, 28'b0000000000000000000000110111, 28'b1111111111111111011100110100, 28'b1111111111111111110111100000, 28'b0000000000000000000000000010, 28'b0000000000000000000101000001, 28'b0000000000000000000000000011, 28'b0000000000000000011100110001, 28'b0000000000000000000000000100, 28'b1111111111111111111101101110, 28'b0000000000000001010100010010, 28'b0000000000000001100000011000, 28'b1111111111111111000111011100, 28'b1111111111111111011011101000, 28'b0000000000000000111111111000, 28'b1111111111111110110001110000, 28'b0000000000000000000111100000, 28'b1111111111111111111111110110, 28'b1111111111111111111111111110, 28'b1111111111111111111111111100, 28'b0000000000000000101111001001}, 
{28'b1111111111111111100010111100, 28'b1111111111111111111111110110, 28'b1111111111111111000010110000, 28'b1111111111111111001100010010, 28'b1111111111111111111100011110, 28'b1111111111111111011101011110, 28'b0000000000000000000000000001, 28'b0000000000000000010111010100, 28'b1111111111111111000010101001, 28'b1111111111111111101010101011, 28'b1111111111111111110011010011, 28'b0000000000000000000000000100, 28'b0000000000000000000111001001, 28'b1111111111111111111101011110, 28'b1111111111111111110000011000, 28'b0000000000000000011000011110, 28'b0000000000000000111001000011, 28'b0000000000000000100001100101, 28'b1111111111111111011110100001, 28'b0000000000000000001100011111, 28'b1111111111111111111100111111, 28'b1111111111111111111000101100, 28'b0000000000000000000101110001, 28'b0000000000000000000100000100, 28'b1111111111111111101110001110, 28'b0000000000000000010110110011, 28'b1111111111111111101000110010, 28'b0000000000000000001111010100, 28'b1111111111111111111111111100, 28'b1111111111111110110100011010, 28'b1111111111111111111001010000, 28'b0000000000000000111001100100}, 
{28'b1111111111111111111001000111, 28'b1111111111111111101010110100, 28'b0000000000000000010011101100, 28'b0000000000000001000000110011, 28'b0000000000000000010101101101, 28'b0000000000000000010101000101, 28'b0000000000000000001011111100, 28'b1111111111111111001100011011, 28'b1111111111111111001011011110, 28'b0000000000000000010001100001, 28'b0000000000000000000011000110, 28'b0000000000000000001011000011, 28'b0000000000000000000101101101, 28'b0000000000000000000001011001, 28'b0000000000000000110100100001, 28'b0000000000000000000001111000, 28'b1111111111111111110010001100, 28'b0000000000000000011010011101, 28'b1111111111111111111000011010, 28'b1111111111111111110110110110, 28'b0000000000000000011100001011, 28'b1111111111111111100000010001, 28'b1111111111111111111001001011, 28'b0000000000000000100000100000, 28'b0000000000000000000101101011, 28'b1111111111111111100100101100, 28'b1111111111111111001101010110, 28'b1111111111111111111100111111, 28'b1111111111111110111000100010, 28'b0000000000000000001111011000, 28'b0000000000000000011010000010, 28'b0000000000000000000000010011}, 
{28'b1111111111111111111100100001, 28'b1111111111111111111010111100, 28'b1111111111111111111100111101, 28'b1111111111111111110111001000, 28'b1111111111111111011110010100, 28'b1111111111111111011100000101, 28'b0000000000000000010000001010, 28'b0000000000000000000010000111, 28'b1111111111111111010001010010, 28'b0000000000000000101010110110, 28'b1111111111111111111010101011, 28'b1111111111111111111111110110, 28'b1111111111111111100011110011, 28'b0000000000000000000001010101, 28'b0000000000000000000111100011, 28'b1111111111111111110010100010, 28'b1111111111111111111011111011, 28'b1111111111111111110101010100, 28'b1111111111111111101011011011, 28'b0000000000000000000000000100, 28'b1111111111111111011100000011, 28'b0000000000000000011010000101, 28'b1111111111111111001001110111, 28'b0000000000000000000001010001, 28'b0000000000000000001010101111, 28'b0000000000000000011111101110, 28'b0000000000000000000110110011, 28'b0000000000000000000001100010, 28'b0000000000000001001010110000, 28'b0000000000000000001101001101, 28'b0000000000000000000000000100, 28'b0000000000000000010101011101}, 
{28'b1111111111111111111011000010, 28'b0000000000000001000000101101, 28'b1111111111111111111111111110, 28'b1111111111111111110111100100, 28'b1111111111111111001001010010, 28'b1111111111111111101100110001, 28'b0000000000000001101001010100, 28'b1111111111111101001111100101, 28'b1111111111111110100110100000, 28'b1111111111111111001100111010, 28'b1111111111111111000111110100, 28'b1111111111111110111111000110, 28'b1111111111111111111111110110, 28'b0000000000000001111011111110, 28'b1111111111111111111001010011, 28'b0000000000000000000000000001, 28'b1111111111111111001001111100, 28'b0000000000000001110010000110, 28'b1111111111111110010110010101, 28'b0000000000000000000000000010, 28'b1111111111111111111111111011, 28'b1111111111111110101001111011, 28'b0000000000000000000000000010, 28'b1111111111111111111111111111, 28'b0000000000000000001110011000, 28'b1111111111111111110001010011, 28'b1111111111111111011010001011, 28'b1111111111111111111111111111, 28'b0000000000000000101100101100, 28'b0000000000000000000000110111, 28'b1111111111111111101011011101, 28'b0000000000000000000000001101}, 
{28'b0000000000000001011110001100, 28'b1111111111111111100011010111, 28'b0000000000000000100001110001, 28'b1111111111111111110111101110, 28'b0000000000000000010011100001, 28'b1111111111111111111111000011, 28'b1111111111111111111111010001, 28'b1111111111111111101000001101, 28'b0000000000000000000000000100, 28'b0000000000000000010111100110, 28'b1111111111111111111111111111, 28'b1111111111111111110000111110, 28'b1111111111111111111111111000, 28'b0000000000000000111010100010, 28'b0000000000000000000100111011, 28'b0000000000000000001010010110, 28'b0000000000000000000110001000, 28'b1111111111111111111001110111, 28'b0000000000000000000101001100, 28'b0000000000000000000000000011, 28'b1111111111111111111101101100, 28'b1111111111111111111111111111, 28'b1111111111111110110001110000, 28'b1111111111111111111111111110, 28'b0000000000000000001110110011, 28'b1111111111111111100010001111, 28'b1111111111111111011101011001, 28'b1111111111111111111111111111, 28'b1111111111111111111111110010, 28'b0000000000000010001110110010, 28'b1111111111111110110110110111, 28'b1111111111111111100010010001}, 
{28'b1111111111111111110100101110, 28'b1111111111111111100101100100, 28'b1111111111111111101111011111, 28'b0000000000000000001001010010, 28'b0000000000000000100011101101, 28'b1111111111111111011110110000, 28'b1111111111111111111111101010, 28'b1111111111111111000111101110, 28'b0000000000000000001111100011, 28'b0000000000000000100010110100, 28'b1111111111111111001001010111, 28'b1111111111111110111111010010, 28'b0000000000000000000110000110, 28'b1111111111111101010001000011, 28'b1111111111111111101100101101, 28'b1111111111111111100000011000, 28'b1111111111111111001101010111, 28'b1111111111111111111111111010, 28'b0000000000000000100010010111, 28'b0000000000000000000000000000, 28'b1111111111111111110100010100, 28'b1111111111111111110100100101, 28'b0000000000000000000000000000, 28'b0000000000000000000000000001, 28'b1111111111111111110000111001, 28'b1111111111111100111110111001, 28'b1111111111111101110001110101, 28'b1111111111111110111010001111, 28'b0000000000000000001110010100, 28'b0000000000000000110100110011, 28'b1111111111111111111111111011, 28'b0000000000000000111101100001}, 
{28'b1111111111111111101000011010, 28'b1111111111111111001001000000, 28'b0000000000000000101001111010, 28'b0000000000000000010011000110, 28'b0000000000000000001011000111, 28'b1111111111111111101000011101, 28'b1111111111111111110111101001, 28'b0000000000000000011001001111, 28'b0000000000000010001001111111, 28'b1111111111111111010100001010, 28'b1111111111111111111111111110, 28'b1111111111111111111111111111, 28'b0000000000000000011110000110, 28'b1111111111111111110001111100, 28'b1111111111111111111011011011, 28'b1111111111111111111011101110, 28'b1111111111111111100110011011, 28'b1111111111111111111111110001, 28'b0000000000000000000000000000, 28'b0000000000000000111010000001, 28'b1111111111111111011101111101, 28'b1111111111111111111111001111, 28'b0000000000000000100000111011, 28'b1111111111111111111101011001, 28'b0000000000000000000000000001, 28'b0000000000000010000110101111, 28'b0000000000000001010011000000, 28'b0000000000000000000000110100, 28'b0000000000000000000000000101, 28'b1111111111111110010100010001, 28'b1111111111111111101110100001, 28'b1111111111111111111111111111}, 
{28'b0000000000000000000011110110, 28'b0000000000000000001100010111, 28'b1111111111111111111100011110, 28'b0000000000000000000000000001, 28'b0000000000000000111011001111, 28'b1111111111111110000100010011, 28'b0000000000000000000000000010, 28'b1111111111111111100111101010, 28'b0000000000000000101111101111, 28'b0000000000000000000000000001, 28'b1111111111111111111011010001, 28'b0000000000000000000000000001, 28'b0000000000000000000000000101, 28'b1111111111111111111111111100, 28'b0000000000000000000001011111, 28'b1111111111111111100100011111, 28'b0000000000000001000010011011, 28'b1111111111111111111110100110, 28'b1111111111111111111100000011, 28'b1111111111111111111111111111, 28'b0000000000000000000000000101, 28'b1111111111111111111110000011, 28'b0000000000000000000000000100, 28'b1111111111111111111111111111, 28'b0000000000000000000011010010, 28'b1111111111111110101110110111, 28'b0000000000000000001101001110, 28'b0000000000000000101110111010, 28'b1111111111111111111111001011, 28'b0000000000000000011000001000, 28'b1111111111111111111111111010, 28'b0000000000000000010011001001}, 
{28'b1111111111111111001100011111, 28'b0000000000000000000010010101, 28'b1111111111111110000100100000, 28'b0000000000000000000001110001, 28'b1111111111111111110011001101, 28'b1111111111111111110101110100, 28'b1111111111111111111111101011, 28'b1111111111111111101000101011, 28'b1111111111111111110110110011, 28'b1111111111111111101111010001, 28'b0000000000000000001100000010, 28'b0000000000000000000110111000, 28'b1111111111111111010010100111, 28'b0000000000000000000000001000, 28'b1111111111111111111111100001, 28'b1111111111111111111101111011, 28'b0000000000000000010010000010, 28'b1111111111111111111010110100, 28'b1111111111111111111000111100, 28'b1111111111111111111000100100, 28'b1111111111111111111111110011, 28'b0000000000000001000101011000, 28'b1111111111111111111111111111, 28'b0000000000000000000000000001, 28'b1111111111111111111101100110, 28'b0000000000000001010001001110, 28'b0000000000000000110000010011, 28'b0000000000000000001000101101, 28'b1111111111111111100111010100, 28'b1111111111111111111101011101, 28'b0000000000000000010000101100, 28'b0000000000000000001110101111}, 
{28'b0000000000000000001000101110, 28'b0000000000000000001010000000, 28'b1111111111111111111111111101, 28'b0000000000000000000000000110, 28'b1111111111111110001000000001, 28'b0000000000000000001011001011, 28'b0000000000000000000110010111, 28'b1111111111111111111111111011, 28'b0000000000000000000000001011, 28'b1111111111111111010100100111, 28'b1111111111111111111111111111, 28'b0000000000000000000000000000, 28'b1111111111111111010110110101, 28'b0000000000000000000000000011, 28'b0000000000000000000000000101, 28'b0000000000000000000000000101, 28'b0000000000000000000000000000, 28'b1111111111111110100100111010, 28'b0000000000000000000010011100, 28'b1111111111111111111111110111, 28'b1111111111111111111111111001, 28'b0000000000000000000000000010, 28'b0000000000000000100001000000, 28'b1111111111111111111111111110, 28'b0000000000000000000000000010, 28'b0000000000000001110100101101, 28'b0000000000000001010111000101, 28'b0000000000000000000000000010, 28'b0000000000000000000000000010, 28'b1111111111111111000100001101, 28'b0000000000000000000000000110, 28'b1111111111111111111111111110}, 
{28'b0000000000000000010011011001, 28'b0000000000000000001101100000, 28'b0000000000000001000000110011, 28'b1111111111111111000000011100, 28'b0000000000000000100001111000, 28'b0000000000000000011110011001, 28'b0000000000000000000001100110, 28'b0000000000000000110001000110, 28'b0000000000000000000011000011, 28'b1111111111111111111100111011, 28'b0000000000000000001001100011, 28'b0000000000000000000001011110, 28'b1111111111111111111111110111, 28'b0000000000000000011110111000, 28'b1111111111111111111110100100, 28'b1111111111111111110101110111, 28'b0000000000000000000000001011, 28'b0000000000000000001000001001, 28'b1111111111111111110011101010, 28'b0000000000000000011001010001, 28'b0000000000000000001000010100, 28'b1111111111111101101011011010, 28'b1111111111111111100010101101, 28'b0000000000000000010111011000, 28'b1111111111111111111111111111, 28'b1111111111111101111110101111, 28'b1111111111111111011111101101, 28'b1111111111111111111010000110, 28'b1111111111111111111111110101, 28'b1111111111111111110001011000, 28'b0000000000000000000000000000, 28'b1111111111111111110101110111}, 
{28'b0000000000000000000000011110, 28'b1111111111111111111111111110, 28'b1111111111111111101000100101, 28'b1111111111111111010100111011, 28'b0000000000000000001010101111, 28'b0000000000000000000000000011, 28'b0000000000000000011000011001, 28'b1111111111111111111110100010, 28'b0000000000000000111111111001, 28'b1111111111111111111110111110, 28'b0000000000000000000000000001, 28'b1111111111111110101000000101, 28'b1111111111111111111111111001, 28'b0000000000000000100000001111, 28'b1111111111111111111111111100, 28'b1111111111111110111101010001, 28'b0000000000000000000000000000, 28'b1111111111111111111101000110, 28'b0000000000000001000011010011, 28'b1111111111111111111111111111, 28'b1111111111111110010000001111, 28'b1111111111111111111111111110, 28'b0000000000000001000010000011, 28'b1111111111111111111111111110, 28'b1111111111111111111111111110, 28'b0000000000000000100011100011, 28'b1111111111111111100111111110, 28'b0000000000000000010001101101, 28'b0000000000000000000000000011, 28'b1111111111111111001100011011, 28'b0000000000000000000000000001, 28'b0000000000000000000000101000}, 
{28'b1111111111111111001000101001, 28'b0000000000000000000000010010, 28'b0000000000000000000000001000, 28'b1111111111111111111110011101, 28'b0000000000000001111110111010, 28'b1111111111111111100000001101, 28'b1111111111111111111110100100, 28'b1111111111111111111110001000, 28'b1111111111111111110100100011, 28'b1111111111111111110011000110, 28'b0000000000000000010000101100, 28'b0000000000000000100010000000, 28'b1111111111111111110110100101, 28'b0000000000000000111111111000, 28'b0000000000000000000000000010, 28'b1111111111111111111111111001, 28'b1111111111111110110111010001, 28'b1111111111111111111111110110, 28'b0000000000000000000000000111, 28'b1111111111111111101011100111, 28'b0000000000000000000000100010, 28'b0000000000000000001001100011, 28'b0000000000000000000011011011, 28'b1111111111111111111101101010, 28'b1111111111111111110010111111, 28'b1111111111111111001100000100, 28'b1111111111111110110100010001, 28'b0000000000000000000000000100, 28'b1111111111111111100011000000, 28'b0000000000000000001010001100, 28'b1111111111111111111111111010, 28'b0000000000000000010011010111}, 
{28'b1111111111111110010110001110, 28'b1111111111111111010111111101, 28'b1111111111111111011000000001, 28'b0000000000000000000000000001, 28'b0000000000000010010010001111, 28'b1111111111111111000111000001, 28'b0000000000000000000000000001, 28'b1111111111111111110010001000, 28'b1111111111111110010111000101, 28'b0000000000000000100011011101, 28'b1111111111111111111111111111, 28'b0000000000000010010001001100, 28'b0000000000000000000000000111, 28'b1111111111111111110011110111, 28'b1111111111111111111111111011, 28'b0000000000000000001000000111, 28'b1111111111111111111011001111, 28'b0000000000000000000000000111, 28'b1111111111111111110100000101, 28'b0000000000000001111110110100, 28'b0000000000000000001001111011, 28'b1111111111111111110101010100, 28'b0000000000000000011100000010, 28'b1111111111111111111111111011, 28'b1111111111111111111111111111, 28'b1111111111111111100111000111, 28'b1111111111111111110100000000, 28'b1111111111111110001000001110, 28'b1111111111111111011011000010, 28'b1111111111111111111111111111, 28'b1111111111111111111111101111, 28'b1111111111111111110000111111}, 
{28'b0000000000000000111001110101, 28'b1111111111111100110011010100, 28'b1111111111111101000110100011, 28'b1111111111111111010100011100, 28'b0000000000000010101011010110, 28'b1111111111111111111111111111, 28'b1111111111111110100111010000, 28'b0000000000000001000011110011, 28'b0000000000000000001111001100, 28'b0000000000000000000000001110, 28'b0000000000000000110101010111, 28'b1111111111111110111010100001, 28'b0000000000000000000000001110, 28'b0000000000000000000001000110, 28'b1111111111111111110111111111, 28'b0000000000000000000100100111, 28'b1111111111111111100101011011, 28'b1111111111111100010100000110, 28'b0000000000000000101010111101, 28'b0000000000000001011000010010, 28'b0000000000000001000011110111, 28'b0000000000000000000000101011, 28'b0000000000000000000111011100, 28'b1111111111111110011000110111, 28'b1111111111111101011110000001, 28'b1111111111111111111110101111, 28'b1111111111111110110011010000, 28'b1111111111111110001010110010, 28'b1111111111111111001110000110, 28'b1111111111111100011111011110, 28'b0000000000000001101011010100, 28'b0000000000000001101101111001}, 
{28'b0000000000000000000000000100, 28'b0000000000000000000000001010, 28'b0000000000000000000000100100, 28'b0000000000000000000000000011, 28'b0000000000000001000010010010, 28'b1111111111111111010000001000, 28'b0000000000000000000100100011, 28'b0000000000000000010010101011, 28'b1111111111111110100110101010, 28'b0000000000000000001001011001, 28'b1111111111111111111110110110, 28'b1111111111111111111111110000, 28'b1111111111111111111111111101, 28'b0000000000000000111101010101, 28'b0000000000000000001101010010, 28'b0000000000000000000101100100, 28'b0000000000000000001111110100, 28'b0000000000000001010101010100, 28'b1111111111111111001000000100, 28'b0000000000000000000000000001, 28'b1111111111111111010101111100, 28'b1111111111111111111111111011, 28'b0000000000000001010000100011, 28'b0000000000000000000010000101, 28'b1111111111111111111111010001, 28'b1111111111111101110000010111, 28'b1111111111111111111101101001, 28'b1111111111111111011000011111, 28'b1111111111111111110000011001, 28'b0000000000000000000000111010, 28'b0000000000000000100010100101, 28'b0000000000000000011010100010}, 
{28'b1111111111111111110100111011, 28'b0000000000000000100010010010, 28'b1111111111111110110010001110, 28'b0000000000000000000101010010, 28'b0000000000000000110001100100, 28'b1111111111111111110101111000, 28'b1111111111111111111110110100, 28'b0000000000000000101001110011, 28'b0000000000000000000000000100, 28'b1111111111111111111111111100, 28'b1111111111111111101111010000, 28'b0000000000000000000000000000, 28'b0000000000000000000000000110, 28'b1111111111111111110111001111, 28'b1111111111111111100000110110, 28'b1111111111111111101111000001, 28'b1111111111111111110001100100, 28'b1111111111111111101111111010, 28'b1111111111111111100011111001, 28'b0000000000000000000000000001, 28'b1111111111111111111111111011, 28'b1111111111111111110100100011, 28'b1111111111111111101110111100, 28'b0000000000000001100101110101, 28'b0000000000000000000000000000, 28'b1111111111111110100011110110, 28'b1111111111111111111101110101, 28'b0000000000000000011111100010, 28'b0000000000000000000000000111, 28'b0000000000000000000000000000, 28'b0000000000000001000000001111, 28'b1111111111111111111111111001}, 
{28'b1111111111111111111111111110, 28'b0000000000000000000001000011, 28'b1111111111111111111111111010, 28'b1111111111111111011000000000, 28'b1111111111111100100011110000, 28'b0000000000000000000000001111, 28'b0000000000000000000000000101, 28'b1111111111111111111110010101, 28'b1111111111111101100110100001, 28'b0000000000000000010100111000, 28'b1111111111111111100110111001, 28'b1111111111111111111111111111, 28'b0000000000000000000000000111, 28'b1111111111111110100001010010, 28'b1111111111111111110100010001, 28'b1111111111111111111111111011, 28'b0000000000000000000000010110, 28'b0000000000000000000010000111, 28'b0000000000000000001001010010, 28'b0000000000000001011000011000, 28'b1111111111111111100001011000, 28'b1111111111111110110011011100, 28'b0000000000000000000000000001, 28'b1111111111111110111101111111, 28'b1111111111111111100110101111, 28'b1111111111111111000100110001, 28'b1111111111111111111110000110, 28'b1111111111111111111100110011, 28'b1111111111111111111011010110, 28'b1111111111111110000111011001, 28'b1111111111111111110111010001, 28'b0000000000000000111110000001}, 
{28'b0000000000000000011100111111, 28'b0000000000000000111000000111, 28'b1111111111111111111111011111, 28'b0000000000000000101000110010, 28'b1111111111111111001010000000, 28'b1111111111111111100000001000, 28'b0000000000000000011000011110, 28'b0000000000000000010001100101, 28'b1111111111111111110011111101, 28'b1111111111111111111111111110, 28'b1111111111111111111111111110, 28'b1111111111111111111111111100, 28'b1111111111111111111111111011, 28'b1111111111111110101101111111, 28'b1111111111111111111111111110, 28'b0000000000000000100100111011, 28'b1111111111111111100010101110, 28'b0000000000000000001000111010, 28'b1111111111111111111111101010, 28'b1111111111111111111111101111, 28'b0000000000000000110101000110, 28'b1111111111111110101100010000, 28'b0000000000000001000111111001, 28'b0000000000000000001100001010, 28'b0000000000000000000000000100, 28'b0000000000000000110110001111, 28'b0000000000000000000000110011, 28'b1111111111111111110110110000, 28'b1111111111111110011110100101, 28'b1111111111111111100011111111, 28'b1111111111111111010100011010, 28'b0000000000000000101101011101}, 
{28'b0000000000000000000000000000, 28'b0000000000000000000001110110, 28'b1111111111111110100010010101, 28'b1111111111111111111111011000, 28'b0000000000000000110100111010, 28'b1111111111111111011011110000, 28'b1111111111111111111100111010, 28'b1111111111111111111111111110, 28'b0000000000000000000101001101, 28'b0000000000000000000000000000, 28'b0000000000000000000000000000, 28'b1111111111111111001011110101, 28'b0000000000000000011000100101, 28'b0000000000000000000001100011, 28'b0000000000000000000000000010, 28'b0000000000000000001001100101, 28'b1111111111111111111111111010, 28'b1111111111111111011001111011, 28'b0000000000000000000100100101, 28'b0000000000000000000000000010, 28'b1111111111111111110111001101, 28'b1111111111111111111010011000, 28'b0000000000000001001011110110, 28'b1111111111111111111111111110, 28'b0000000000000000000000000001, 28'b1111111111111110110101000101, 28'b1111111111111110101100010100, 28'b0000000000000000111101110011, 28'b1111111111111111111111101011, 28'b1111111111111111111111111010, 28'b0000000000000000000111000101, 28'b0000000000000001001000010110}, 
{28'b1111111111111110101000110001, 28'b1111111111111111111111111111, 28'b1111111111111111001001100011, 28'b0000000000000000000001000110, 28'b1111111111111110100101100010, 28'b0000000000000000000000000000, 28'b1111111111111111111111111011, 28'b1111111111111111101111010001, 28'b1111111111111101110111101110, 28'b1111111111111111111001011010, 28'b0000000000000000000000000001, 28'b1111111111111111111101111000, 28'b1111111111111111111111111010, 28'b0000000000000000000000000001, 28'b1111111111111111111101110011, 28'b1111111111111111110011010001, 28'b1111111111111111011010001111, 28'b1111111111111111100111100101, 28'b0000000000000000010000111100, 28'b1111111111111111111111011000, 28'b1111111111111111111001100001, 28'b0000000000000000000000000001, 28'b0000000000000001010110001100, 28'b1111111111111111111111111101, 28'b0000000000000000100110010000, 28'b0000000000000000010111011110, 28'b1111111111111111011100110001, 28'b0000000000000000110110100110, 28'b1111111111111111110100010010, 28'b0000000000000000000000000000, 28'b1111111111111111111111101101, 28'b0000000000000010010101000000}, 
{28'b1111111111111110101111100111, 28'b0000000000000000000111100110, 28'b0000000000000000001100111110, 28'b1111111111111111111000110100, 28'b0000000000000000111110100001, 28'b1111111111111110110010101000, 28'b1111111111111111111110001101, 28'b0000000000000001000011111111, 28'b0000000000000000101000110010, 28'b0000000000000000000010010110, 28'b1111111111111111111111111110, 28'b1111111111111111101110011110, 28'b1111111111111111101001000110, 28'b1111111111111111101111011100, 28'b1111111111111111110011010010, 28'b0000000000000000010111000110, 28'b1111111111111111111111111110, 28'b0000000000000000000010000100, 28'b0000000000000000100100001011, 28'b0000000000000000000000000001, 28'b0000000000000000000000000001, 28'b0000000000000000000011110100, 28'b0000000000000001000000100000, 28'b0000000000000000001011101101, 28'b0000000000000000000001101101, 28'b1111111111111111100100011101, 28'b1111111111111111111111111110, 28'b0000000000000000000000000000, 28'b1111111111111111111100011000, 28'b1111111111111111111100111010, 28'b1111111111111111111111111011, 28'b0000000000000000010001010011}, 
{28'b1111111111111111111111111101, 28'b0000000000000000000000111111, 28'b1111111111111111001001101110, 28'b1111111111111111101100111011, 28'b0000000000000001001000001110, 28'b1111111111111111111111111010, 28'b1111111111111111101100001011, 28'b0000000000000000111110100101, 28'b1111111111111111110010011100, 28'b0000000000000001001010101010, 28'b0000000000000000010101111001, 28'b1111111111111111100001001110, 28'b0000000000000000000000001001, 28'b0000000000000000000000111001, 28'b1111111111111111111100001111, 28'b0000000000000000000101011100, 28'b1111111111111111101100010001, 28'b1111111111111110111100100110, 28'b0000000000000001000111001001, 28'b0000000000000000100111110001, 28'b0000000000000010100010011111, 28'b0000000000000000110011011000, 28'b0000000000000000111111100000, 28'b1111111111111111111111111100, 28'b0000000000000000000000000000, 28'b0000000000000000000000000000, 28'b0000000000000000001110101011, 28'b0000000000000000010100010010, 28'b1111111111111110010100011111, 28'b1111111111111111111111111100, 28'b1111111111111111111110101100, 28'b1111111111111111111110010100}, 
{28'b0000000000000000000000001000, 28'b1111111111111111101001100100, 28'b1111111111111111100101011111, 28'b0000000000000000000000000000, 28'b1111111111111111000001101000, 28'b0000000000000000000000000001, 28'b0000000000000000110001000000, 28'b0000000000000000011011111100, 28'b0000000000000000001101100110, 28'b1111111111111111100110101110, 28'b0000000000000000000000000001, 28'b1111111111111111111111111111, 28'b1111111111111111111111111100, 28'b1111111111111111111111111101, 28'b1111111111111111110101000101, 28'b0000000000000000110011101110, 28'b1111111111111111111111111111, 28'b1111111111111111111111110111, 28'b1111111111111110110010100110, 28'b0000000000000000000000000010, 28'b1111111111111111001110101111, 28'b1111111111111111111111101111, 28'b0000000000000000000000000010, 28'b1111111111111111111110111100, 28'b0000000000000000000011110111, 28'b0000000000000000000100011101, 28'b0000000000000000000111001001, 28'b0000000000000000100011011011, 28'b1111111111111111101111010111, 28'b1111111111111111111110000010, 28'b1111111111111110001101001001, 28'b0000000000000000010100001011}, 
{28'b0000000000000001110001000110, 28'b1111111111111111111101110001, 28'b0000000000000000010000111101, 28'b1111111111111111100101001100, 28'b1111111111111111101010001001, 28'b0000000000000000001000100010, 28'b0000000000000000101001000001, 28'b0000000000000000000000000001, 28'b0000000000000010000110111010, 28'b0000000000000000000000000101, 28'b1111111111111111111010100001, 28'b0000000000000000000100110101, 28'b0000000000000000011000000101, 28'b1111111111111111111111010101, 28'b0000000000000000001101101000, 28'b0000000000000000011010011100, 28'b1111111111111111111110111001, 28'b1111111111111110001110000010, 28'b1111111111111111110001100100, 28'b1111111111111111111111100100, 28'b0000000000000000011101110001, 28'b0000000000000000000000011011, 28'b1111111111111111111111111000, 28'b0000000000000000011100110011, 28'b0000000000000000000100100110, 28'b1111111111111110111100100001, 28'b1111111111111111100101101101, 28'b0000000000000000100001110110, 28'b1111111111111111111000110001, 28'b0000000000000001000010000100, 28'b1111111111111111111111101110, 28'b1111111111111111010010001111}, 
{28'b0000000000000000000011010100, 28'b0000000000000000011010000101, 28'b1111111111111111111111111111, 28'b1111111111111111110110000101, 28'b1111111111111110100101101001, 28'b1111111111111111111111111001, 28'b0000000000000000001011110010, 28'b1111111111111111110100001101, 28'b0000000000000000101010001101, 28'b1111111111111111110111010000, 28'b1111111111111111111111110010, 28'b1111111111111111110111011100, 28'b1111111111111111111111111100, 28'b1111111111111111110110100001, 28'b0000000000000000000000000001, 28'b0000000000000001010000001001, 28'b0000000000000000000000000001, 28'b1111111111111111111111100011, 28'b1111111111111111111111111100, 28'b1111111111111111111111111101, 28'b1111111111111111111111111100, 28'b1111111111111111111111111001, 28'b0000000000000000001000101110, 28'b0000000000000000100000001110, 28'b0000000000000000000000000000, 28'b0000000000000000000001000100, 28'b0000000000000000001000010010, 28'b1111111111111111111111110111, 28'b0000000000000000000000000001, 28'b0000000000000000000101001110, 28'b0000000000000000000000011000, 28'b0000000000000000011000110010}, 
{28'b1111111111111110110000111100, 28'b0000000000000000100001010110, 28'b0000000000000000000100100110, 28'b1111111111111111100101000111, 28'b1111111111111110011001110010, 28'b1111111111111111111011010100, 28'b0000000000000000010001001001, 28'b1111111111111110011010010000, 28'b0000000000000010000010111101, 28'b0000000000000000010010010110, 28'b0000000000000000000100000000, 28'b0000000000000000011000001000, 28'b0000000000000000001011010110, 28'b0000000000000000000000001011, 28'b0000000000000001101000011001, 28'b1111111111111111101010011101, 28'b0000000000000000000001010101, 28'b0000000000000000000000000001, 28'b1111111111111111111110010010, 28'b0000000000000000000000111101, 28'b1111111111111110010001011110, 28'b0000000000000000000100010101, 28'b0000000000000000100111001001, 28'b0000000000000000001001100111, 28'b0000000000000000001001001111, 28'b1111111111111101010111111111, 28'b1111111111111110101000101111, 28'b1111111111111111000010011001, 28'b0000000000000000000000101011, 28'b1111111111111111111111100011, 28'b0000000000000001010011011011, 28'b1111111111111111001011100101}, 
{28'b1111111111111111111100101101, 28'b1111111111111111001110001111, 28'b1111111111111111100101100010, 28'b1111111111111110010111011000, 28'b1111111111111110111101011001, 28'b0000000000000001010110000100, 28'b0000000000000001001111010101, 28'b1111111111111111010100011101, 28'b0000000000000000001010101001, 28'b1111111111111111110110000100, 28'b1111111111111111100111111101, 28'b1111111111111110111111101001, 28'b0000000000000000011010011001, 28'b1111111111111110110111010000, 28'b0000000000000000110000010100, 28'b1111111111111111111111111010, 28'b0000000000000001010101111111, 28'b1111111111111111111111111111, 28'b1111111111111111111110000000, 28'b1111111111111111011101010110, 28'b1111111111111111110101010110, 28'b1111111111111111101111011111, 28'b1111111111111110111011111111, 28'b0000000000000000010101000101, 28'b1111111111111111111111111110, 28'b1111111111111111111110011000, 28'b1111111111111111000101100101, 28'b0000000000000001010000100110, 28'b0000000000000001000111011100, 28'b1111111111111111101000110110, 28'b1111111111111101011110100101, 28'b0000000000000000100100100100}, 
{28'b0000000000000000000000000110, 28'b1111111111111111111001011101, 28'b1111111111111111111111111100, 28'b1111111111111111100111000111, 28'b0000000000000000000111010010, 28'b0000000000000000000010010101, 28'b0000000000000000010001110101, 28'b0000000000000000000001011110, 28'b0000000000000000011110001011, 28'b1111111111111111111111110000, 28'b0000000000000000000000000000, 28'b0000000000000000011000011011, 28'b0000000000000000000000011110, 28'b0000000000000000000011001000, 28'b1111111111111111011110000111, 28'b1111111111111111100100011011, 28'b0000000000000000000000000001, 28'b0000000000000000101110100001, 28'b0000000000000000001110100010, 28'b0000000000000000100000001100, 28'b1111111111111111111011110001, 28'b1111111111111111010111000101, 28'b1111111111111111111111111101, 28'b0000000000000000010011000001, 28'b1111111111111111111111111101, 28'b0000000000000000001000010010, 28'b1111111111111111111110110001, 28'b0000000000000000010001010010, 28'b0000000000000000000000000011, 28'b0000000000000000010101010010, 28'b1111111111111110011110110110, 28'b1111111111111111111111111110}, 
{28'b0000000000000001001111011101, 28'b1111111111111111111101101100, 28'b0000000000000000100110011000, 28'b1111111111111110110001110111, 28'b1111111111111111001110100100, 28'b1111111111111111111111111110, 28'b1111111111111111111111111101, 28'b0000000000000000000111000000, 28'b0000000000000000000000100110, 28'b1111111111111111011111110000, 28'b0000000000000000000000000000, 28'b0000000000000000000000100000, 28'b0000000000000000000000000000, 28'b0000000000000000000000000101, 28'b1111111111111111011110111100, 28'b0000000000000000100100100000, 28'b1111111111111111111111100101, 28'b1111111111111111111000000101, 28'b0000000000000000000000000010, 28'b0000000000000000011110101110, 28'b1111111111111111001100100110, 28'b0000000000000000011101101111, 28'b0000000000000000100011110111, 28'b0000000000000000100001000001, 28'b1111111111111111111111111111, 28'b0000000000000010001101001011, 28'b1111111111111111011000110011, 28'b0000000000000001011101000010, 28'b1111111111111111110010110011, 28'b1111111111111110100011101011, 28'b1111111111111111010011100111, 28'b0000000000000000100011101100}, 
{28'b1111111111111101110100111101, 28'b1111111111111111111001001010, 28'b1111111111111111011000100100, 28'b1111111111111111111111111111, 28'b0000000000000001000010110000, 28'b1111111111111111010010010011, 28'b1111111111111111110000101010, 28'b0000000000000000111100111111, 28'b0000000000000000011000001101, 28'b1111111111111111000011000101, 28'b0000000000000000000000000010, 28'b1111111111111111111000110011, 28'b1111111111111111111101011111, 28'b0000000000000000100011001101, 28'b1111111111111111000001000110, 28'b1111111111111111111101001000, 28'b0000000000000000000000000000, 28'b1111111111111111111111110101, 28'b1111111111111111111011111001, 28'b0000000000000000000000000001, 28'b1111111111111111001111010101, 28'b1111111111111111111111111100, 28'b0000000000000000000000000001, 28'b1111111111111110101011111100, 28'b0000000000000000010001111110, 28'b0000000000000010011110101011, 28'b0000000000000001011000100010, 28'b1111111111111111110110110101, 28'b1111111111111111010110111001, 28'b1111111111111110001101001001, 28'b0000000000000000000000000101, 28'b1111111111111111110011100000}, 
{28'b0000000000000000000101011111, 28'b0000000000000000110110101101, 28'b0000000000000000000101011100, 28'b1111111111111111011001010100, 28'b0000000000000000000001001011, 28'b1111111111111111111001011111, 28'b0000000000000000000000000011, 28'b0000000000000000110101010111, 28'b0000000000000000110111000001, 28'b1111111111111111011101110010, 28'b0000000000000000100011111101, 28'b0000000000000000000110001001, 28'b1111111111111111111111111110, 28'b1111111111111111111100010110, 28'b1111111111111111010111010110, 28'b0000000000000001000000110000, 28'b1111111111111111110101001001, 28'b1111111111111110101101010010, 28'b0000000000000000011101010001, 28'b1111111111111111111111111101, 28'b1111111111111111111111111100, 28'b0000000000000000011101111010, 28'b1111111111111111101100111110, 28'b1111111111111111111110110001, 28'b1111111111111111110010110010, 28'b0000000000000000010110100100, 28'b1111111111111111011100000101, 28'b0000000000000000100010010101, 28'b1111111111111110100010111000, 28'b0000000000000000010100100110, 28'b1111111111111111111111111000, 28'b0000000000000000101000000110}, 
{28'b1111111111111111110101000001, 28'b0000000000000000000000001001, 28'b0000000000000000010110110010, 28'b0000000000000000000000000001, 28'b1111111111111111110000011000, 28'b1111111111111111111111010001, 28'b0000000000000000011010010001, 28'b1111111111111111111111111111, 28'b0000000000000000000000000011, 28'b0000000000000000000001010011, 28'b0000000000000000000000000010, 28'b0000000000000000000101000110, 28'b1111111111111111100100110010, 28'b0000000000000000000010101010, 28'b0000000000000000011100010110, 28'b0000000000000000001011111101, 28'b0000000000000000011011000001, 28'b1111111111111111111111110111, 28'b1111111111111111111111101010, 28'b0000000000000000100000110001, 28'b0000000000000000111111010101, 28'b1111111111111111100110111101, 28'b0000000000000000000000000001, 28'b1111111111111111111111011110, 28'b0000000000000000000010111011, 28'b1111111111111110001001111111, 28'b1111111111111111111111110010, 28'b1111111111111111101101111000, 28'b1111111111111111111111111100, 28'b0000000000000010010000100010, 28'b0000000000000000000000000100, 28'b1111111111111111001011010010}, 
{28'b1111111111111111111001001000, 28'b1111111111111111100001011100, 28'b1111111111111111111101101111, 28'b0000000000000000000001110010, 28'b0000000000000000010111001110, 28'b1111111111111111111111111110, 28'b0000000000000000000000000011, 28'b1111111111111111111010000100, 28'b0000000000000000010010000101, 28'b1111111111111111111101111001, 28'b0000000000000000000000000010, 28'b0000000000000000001000000110, 28'b0000000000000001001011100001, 28'b1111111111111111100101111001, 28'b0000000000000000000011001110, 28'b1111111111111100100110110110, 28'b1111111111111111111101001001, 28'b1111111111111111110000100001, 28'b0000000000000000000010000011, 28'b1111111111111111110011001110, 28'b0000000000000000010111100011, 28'b1111111111111111000110101000, 28'b0000000000000000011101001110, 28'b0000000000000000011010111111, 28'b1111111111111111111100101001, 28'b1111111111111101001001111110, 28'b1111111111111111000101011111, 28'b1111111111111111111010011010, 28'b1111111111111111111011010011, 28'b0000000000000001100011111110, 28'b1111111111111111111110100000, 28'b0000000000000000100111011100}, 
{28'b0000000000000000001100000001, 28'b0000000000000000000000000010, 28'b0000000000000000101100100101, 28'b1111111111111111100010111101, 28'b1111111111111111101110011001, 28'b0000000000000000111100111001, 28'b1111111111111111010111000100, 28'b0000000000000000001110101110, 28'b1111111111111110110000110010, 28'b0000000000000000000010001111, 28'b0000000000000000000100010010, 28'b1111111111111111101010100001, 28'b0000000000000000000000001000, 28'b0000000000000000000000000000, 28'b1111111111111111001111111010, 28'b0000000000000001101110101101, 28'b1111111111111111000000110101, 28'b1111111111111111111100111100, 28'b0000000000000000011110011011, 28'b1111111111111111111111111101, 28'b0000000000000000010001101111, 28'b1111111111111110000101010110, 28'b0000000000000001010000001011, 28'b1111111111111111111111111111, 28'b1111111111111111100000010011, 28'b0000000000000001111100000100, 28'b0000000000000000100101011001, 28'b1111111111111111010111100111, 28'b1111111111111111011101100101, 28'b1111111111111101110110011111, 28'b1111111111111111111101011001, 28'b0000000000000000000100000100}, 
{28'b1111111111111111111111111111, 28'b0000000000000000000001101011, 28'b1111111111111111110111000110, 28'b1111111111111110111011011001, 28'b1111111111111111111111111010, 28'b1111111111111110011011100010, 28'b0000000000000000000000000100, 28'b0000000000000001001101101110, 28'b0000000000000000111110100010, 28'b0000000000000000000100110101, 28'b0000000000000000000000000000, 28'b1111111111111111100011110011, 28'b0000000000000001010101000001, 28'b1111111111111111111111111111, 28'b1111111111111111111111111010, 28'b1111111111111111111111111001, 28'b0000000000000001101111000101, 28'b0000000000000000000000011010, 28'b1111111111111111110101110101, 28'b1111111111111111110010111011, 28'b1111111111111110101101100110, 28'b0000000000000000100001101100, 28'b0000000000000000000000000000, 28'b0000000000000000000000000000, 28'b0000000000000000001000000110, 28'b1111111111111111101101110010, 28'b1111111111111110001010000101, 28'b0000000000000001000110101000, 28'b1111111111111110001110011111, 28'b0000000000000000001101000101, 28'b1111111111111111101011110010, 28'b0000000000000000000000000000}, 
{28'b0000000000000000001111101100, 28'b0000000000000000101111101110, 28'b0000000000000000000010011110, 28'b1111111111111111111111001111, 28'b1111111111111110001010011011, 28'b0000000000000000000000001110, 28'b1111111111111111111111111111, 28'b0000000000000000111110000001, 28'b0000000000000001000110111011, 28'b1111111111111111111111111101, 28'b1111111111111111111111111101, 28'b1111111111111111111111101011, 28'b0000000000000000000000000010, 28'b0000000000000000000000100001, 28'b0000000000000000000000000000, 28'b0000000000000000000000000011, 28'b0000000000000000000000000111, 28'b1111111111111111111111110101, 28'b0000000000000000101011100000, 28'b1111111111111111100101101001, 28'b1111111111111110010001011010, 28'b1111111111111111110111100001, 28'b1111111111111111100110101100, 28'b1111111111111111100111111110, 28'b1111111111111111101110010001, 28'b1111111111111111111111110001, 28'b1111111111111111101111111001, 28'b1111111111111111111010011001, 28'b1111111111111111111101010101, 28'b0000000000000000100100001101, 28'b1111111111111111111111111010, 28'b0000000000000001110110101001}
};

localparam logic signed [27:0] bias [32] = '{
28'b0000000000000101111001011010,  // 1.474280834197998
28'b0000000000000010110001000001,  // 0.6914801001548767
28'b0000000000000101110000110011,  // 1.4406442642211914
28'b0000000000000101101000011101,  // 1.408045768737793
28'b0000000000000011111100100010,  // 0.9864811301231384
28'b0000000000000011011101000101,  // 0.8636202812194824
28'b1111111111111101100010011101,  // -0.6153604388237
28'b0000000000000001111011111000,  // 0.4839226007461548
28'b0000000000000001111100011111,  // 0.4862793982028961
28'b0000000000000001011111001000,  // 0.37162142992019653
28'b0000000000000001110101101110,  // 0.45989668369293213
28'b0000000000000101001100110000,  // 1.2998151779174805
28'b1111111111111011111011110001,  // -1.016528844833374
28'b1111111111111110100101110000,  // -0.35249894857406616
28'b0000000000000001110010001000,  // 0.44582197070121765
28'b1111111111111111100011010101,  // -0.1119980737566948
28'b1111111111111111101110110011,  // -0.06717441976070404
28'b0000000000000000000001001111,  // 0.00487547367811203
28'b0000000000000000110001110101,  // 0.1946917623281479
28'b1111111111111100111000011001,  // -0.7796769738197327
28'b0000000000000010111010100011,  // 0.7287401556968689
28'b0000000000000110110111000000,  // 1.714877724647522
28'b1111111111111001100111001001,  // -1.5971007347106934
28'b0000000000000000010010111011,  // 0.07393483817577362
28'b0000000000000001010010100100,  // 0.3225609362125397
28'b0000000000000011011000011001,  // 0.8453295230865479
28'b0000000000000011100110000010,  // 0.898597240447998
28'b0000000000000001000001001111,  // 0.2548799514770508
28'b0000000000000011111001001110,  // 0.9735668301582336
28'b0000000000000100100000010011,  // 1.1261906623840332
28'b0000000000000001110010100110,  // 0.44768181443214417
28'b1111111111110110100001111001   // -2.3676068782806396
};
endpackage