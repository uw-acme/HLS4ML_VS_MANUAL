// Width: 12
// NFRAC: 6
package dense_2_12_6;

localparam logic signed [11:0] weights [64][32] = '{ 
{12'b000000010001, 12'b000000000000, 12'b111111110011, 12'b111111111110, 12'b000000010000, 12'b000000000000, 12'b111111110110, 12'b111111111111, 12'b111111101110, 12'b000000000101, 12'b000000000000, 12'b111111111111, 12'b111111111111, 12'b111111110011, 12'b111111111100, 12'b111111101111, 12'b000000000000, 12'b111111111111, 12'b111111110011, 12'b111111110101, 12'b000000000000, 12'b000000000000, 12'b111111111111, 12'b111111111111, 12'b000000000000, 12'b000000000110, 12'b000000011000, 12'b000000001011, 12'b111111111111, 12'b000000000011, 12'b111111100101, 12'b000000000000}, 
{12'b111111111001, 12'b111111110110, 12'b111111110111, 12'b111111111100, 12'b111111111111, 12'b000000000010, 12'b111111110001, 12'b000000000000, 12'b000000000000, 12'b111111111011, 12'b000000001001, 12'b111111111101, 12'b111111111100, 12'b111111110010, 12'b000000000000, 12'b111111111100, 12'b000000000000, 12'b111111110011, 12'b000000001010, 12'b000000001110, 12'b111111111101, 12'b111111111111, 12'b111111111111, 12'b000000000001, 12'b111111111011, 12'b000000010001, 12'b000000001111, 12'b000000000000, 12'b000000000001, 12'b111111100000, 12'b000000000000, 12'b000000000000}, 
{12'b000000000100, 12'b111111111000, 12'b111111110111, 12'b111111111101, 12'b111111111011, 12'b111111111010, 12'b111111110100, 12'b000000000000, 12'b111111110111, 12'b000000000000, 12'b000000000000, 12'b111111111010, 12'b000000000101, 12'b111111111011, 12'b111111111111, 12'b111111111101, 12'b000000000000, 12'b000000000110, 12'b000000000011, 12'b000000001110, 12'b000000000010, 12'b111111111010, 12'b000000000000, 12'b000000000010, 12'b111111111110, 12'b000000001101, 12'b000000001001, 12'b000000000110, 12'b111111111111, 12'b111111110110, 12'b111111111111, 12'b000000000110}, 
{12'b000000001000, 12'b000000000001, 12'b000000000011, 12'b111111111111, 12'b111111011111, 12'b000000000000, 12'b000000000000, 12'b000000001110, 12'b000000001111, 12'b111111111111, 12'b111111111111, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b111111111110, 12'b000000001101, 12'b000000000000, 12'b111111111110, 12'b111111111111, 12'b111111110100, 12'b111111111100, 12'b000000000011, 12'b111111111011, 12'b111111111111, 12'b000000000000, 12'b111111111100, 12'b000000000100, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111110010, 12'b000000010011}, 
{12'b111111010100, 12'b111111111110, 12'b111111111111, 12'b000000000000, 12'b111111111110, 12'b000000000000, 12'b111111111100, 12'b111111110110, 12'b000000000011, 12'b111111111110, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b000000001101, 12'b000000000000, 12'b000000010101, 12'b111111111111, 12'b000000001101, 12'b111111100110, 12'b000000000000, 12'b111111111000, 12'b000000001010, 12'b000000010000, 12'b000000000000, 12'b000000000010, 12'b000000001010, 12'b000000001111, 12'b000000000001, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b000000001110}, 
{12'b000000000011, 12'b111111111111, 12'b000000001001, 12'b111111010110, 12'b111110100111, 12'b111111101001, 12'b000000010110, 12'b111111011000, 12'b111111111111, 12'b111111010100, 12'b111111011111, 12'b111111101010, 12'b000000010110, 12'b111111111111, 12'b111111111111, 12'b000000000000, 12'b111111111111, 12'b111111111111, 12'b111111110111, 12'b111111111111, 12'b111111100000, 12'b000000000000, 12'b000000001011, 12'b111111111111, 12'b000000000001, 12'b000000010001, 12'b000000000011, 12'b111111111111, 12'b111111111111, 12'b000000001101, 12'b111111111101, 12'b000000001100}, 
{12'b111111111101, 12'b111111110101, 12'b111111110000, 12'b111111111100, 12'b111111101101, 12'b000000000100, 12'b111111110100, 12'b111111110110, 12'b111111100101, 12'b000000000011, 12'b111111111111, 12'b111111110101, 12'b000000000111, 12'b111111111111, 12'b111111111101, 12'b111111011100, 12'b111111111111, 12'b000000000101, 12'b000000001100, 12'b111111110101, 12'b111111110110, 12'b111111111011, 12'b111111111111, 12'b000000000001, 12'b111111111101, 12'b111111010110, 12'b111111101111, 12'b111111111101, 12'b000000000000, 12'b111111111110, 12'b000000000001, 12'b111111111111}, 
{12'b111111110110, 12'b111111111010, 12'b111111111010, 12'b111111110000, 12'b111111111000, 12'b111111111111, 12'b000000000110, 12'b111111111010, 12'b000000001100, 12'b000000000000, 12'b000000000000, 12'b111111111111, 12'b000000001110, 12'b000000000000, 12'b111111111111, 12'b111111111011, 12'b111111111111, 12'b000000000000, 12'b111111111111, 12'b000000000000, 12'b111111111111, 12'b111111111111, 12'b000000000000, 12'b111111111111, 12'b000000000010, 12'b111111110100, 12'b000000000000, 12'b111111111111, 12'b111111111011, 12'b111111111111, 12'b000000000000, 12'b111111111111}, 
{12'b111111100001, 12'b111111111100, 12'b111111100111, 12'b000000000111, 12'b000000011111, 12'b111111111111, 12'b111111111110, 12'b000000001111, 12'b111111100011, 12'b111111111101, 12'b000000000000, 12'b111111110011, 12'b111111111111, 12'b000000000100, 12'b111111110011, 12'b000000110000, 12'b111111111111, 12'b000000000010, 12'b000000001101, 12'b000000001111, 12'b000000000000, 12'b111111101010, 12'b000000000000, 12'b000000011010, 12'b111111110100, 12'b000000101100, 12'b111111110110, 12'b111111110010, 12'b111111100001, 12'b111111100010, 12'b000000000000, 12'b000000000011}, 
{12'b000000000000, 12'b111111111111, 12'b111111111011, 12'b000000000000, 12'b000000010011, 12'b111111111110, 12'b111111111011, 12'b000000000101, 12'b000000000110, 12'b000000000000, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111000, 12'b111111111111, 12'b000000000000, 12'b000000000000, 12'b111111111111, 12'b000000000000, 12'b000000000101, 12'b000000000001, 12'b111111111111, 12'b000000000000, 12'b000000000000, 12'b000000000010, 12'b111111110111, 12'b000000000100, 12'b000000001111, 12'b111111111111, 12'b000000000000, 12'b000000000011, 12'b000000000100}, 
{12'b000000000110, 12'b000000000000, 12'b111111111001, 12'b111111101111, 12'b111111001101, 12'b000000001000, 12'b000000000000, 12'b111111001011, 12'b000000000010, 12'b111111111111, 12'b000000000000, 12'b111111111111, 12'b000000000000, 12'b000000000000, 12'b111111111110, 12'b111111100111, 12'b111111111111, 12'b000000001110, 12'b000000001000, 12'b000000001100, 12'b111111100011, 12'b111111101001, 12'b000000000111, 12'b111111111101, 12'b111111111101, 12'b000000010110, 12'b111111111001, 12'b111111111111, 12'b111111111111, 12'b000000001101, 12'b111111111111, 12'b000000000000}, 
{12'b111111110011, 12'b111111100000, 12'b000000000000, 12'b111111111111, 12'b000000010101, 12'b111111101110, 12'b111111110001, 12'b000000000111, 12'b111111111111, 12'b000000001001, 12'b000000000100, 12'b111111111011, 12'b000000000000, 12'b000000000000, 12'b111111111110, 12'b111111101111, 12'b000000001011, 12'b000000000001, 12'b000000010011, 12'b000000000101, 12'b000000000000, 12'b111111111101, 12'b000000001000, 12'b111111111010, 12'b111111101100, 12'b111111111111, 12'b000000001011, 12'b111111111111, 12'b000000000000, 12'b111111111001, 12'b000000001000, 12'b000000010001}, 
{12'b000000000000, 12'b000000000000, 12'b000000001110, 12'b000000000000, 12'b111111111101, 12'b000000001011, 12'b000000000101, 12'b111111111111, 12'b000000000000, 12'b111111110111, 12'b111111111100, 12'b111111110101, 12'b111111111111, 12'b000000000011, 12'b111111111011, 12'b000000110101, 12'b000000000000, 12'b111111111001, 12'b111111110011, 12'b111111111111, 12'b000000001100, 12'b000000001000, 12'b000000000000, 12'b111111111111, 12'b000000001110, 12'b000000010001, 12'b000000011111, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b111111111111, 12'b111111111011}, 
{12'b111111110110, 12'b000000000011, 12'b000000000010, 12'b111111110000, 12'b111111101110, 12'b000000011110, 12'b000000000011, 12'b000000000000, 12'b111111110101, 12'b111111111010, 12'b000000001000, 12'b000000000100, 12'b000000000000, 12'b111111111010, 12'b000000010010, 12'b111111111111, 12'b111111111111, 12'b000000000000, 12'b000000000000, 12'b111111111101, 12'b000000000101, 12'b000000000001, 12'b000000000111, 12'b111111111111, 12'b000000000000, 12'b000000101010, 12'b111111111100, 12'b111111111110, 12'b111111111111, 12'b111111111001, 12'b111111111101, 12'b000000001011}, 
{12'b000000000011, 12'b000000000100, 12'b000000010100, 12'b111111111101, 12'b000000000110, 12'b000000010110, 12'b000000000000, 12'b111111111110, 12'b000000000111, 12'b111111111000, 12'b111111111111, 12'b111111111000, 12'b000000000000, 12'b000000011001, 12'b111111111110, 12'b000000000000, 12'b000000001111, 12'b000000000000, 12'b000000000000, 12'b111111101011, 12'b111111110000, 12'b111111111101, 12'b111111111111, 12'b111111110110, 12'b111111111101, 12'b111111111010, 12'b111111110011, 12'b111111110010, 12'b000000000001, 12'b000000000111, 12'b111111100110, 12'b000000000000}, 
{12'b111111101100, 12'b000000000000, 12'b111111111111, 12'b111111111100, 12'b111111111111, 12'b000000001000, 12'b111111111011, 12'b000000010001, 12'b111111101000, 12'b111111111111, 12'b000000000000, 12'b111111111111, 12'b000000000000, 12'b000000000000, 12'b111111111111, 12'b111111111010, 12'b000000000101, 12'b000000001011, 12'b111111111111, 12'b111111101111, 12'b111111111100, 12'b000000000111, 12'b000000000100, 12'b000000000000, 12'b000000000000, 12'b000000000101, 12'b111111110000, 12'b000000000000, 12'b111111111111, 12'b000000000000, 12'b000000000000, 12'b111111110111}, 
{12'b111111101010, 12'b111111111111, 12'b111111111111, 12'b111111111110, 12'b111111111111, 12'b000000000110, 12'b000000000000, 12'b000000000010, 12'b000000000010, 12'b000000000100, 12'b000000000101, 12'b000000001010, 12'b000000000001, 12'b111111111001, 12'b000000000000, 12'b000000011000, 12'b000000000000, 12'b000000000000, 12'b111111111111, 12'b000000000111, 12'b000000001001, 12'b000000000001, 12'b000000000010, 12'b111111111110, 12'b111111111101, 12'b000000000001, 12'b111111111011, 12'b111111110111, 12'b000000001101, 12'b111111111110, 12'b000000000010, 12'b111111110011}, 
{12'b000000000000, 12'b111111111111, 12'b000000000010, 12'b000000000000, 12'b000000111010, 12'b111111111111, 12'b000000000000, 12'b111111111111, 12'b000000000111, 12'b111111111011, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000001000, 12'b000000000000, 12'b111111110110, 12'b111111111111, 12'b111111111011, 12'b000000010100, 12'b000000000000, 12'b111111111111, 12'b111111111111, 12'b000000000000, 12'b111111111111, 12'b000000000000, 12'b000000000100, 12'b000000000000, 12'b000000000000, 12'b111111111111, 12'b111111111111, 12'b000000000000, 12'b000000000010}, 
{12'b111111111111, 12'b000000000001, 12'b111111111111, 12'b000000000011, 12'b111111111101, 12'b111111111000, 12'b111111111100, 12'b000000010001, 12'b000000000000, 12'b000000000110, 12'b111111111111, 12'b000000000100, 12'b111111111101, 12'b111111110101, 12'b111111110011, 12'b000000000000, 12'b111111111111, 12'b111111111101, 12'b000000000000, 12'b000000000000, 12'b111111111111, 12'b000000000100, 12'b000000000010, 12'b111111110111, 12'b000000000111, 12'b111111110101, 12'b000000000000, 12'b000000000000, 12'b111111110101, 12'b000000000000, 12'b000000000010, 12'b111111111110}, 
{12'b111111111111, 12'b111111111001, 12'b000000000000, 12'b111111111100, 12'b000000001101, 12'b111111111111, 12'b111111111110, 12'b000000000110, 12'b111111100110, 12'b000000000000, 12'b111111111101, 12'b111111111111, 12'b000000010110, 12'b000000001110, 12'b111111111001, 12'b111111111110, 12'b111111111111, 12'b000000000000, 12'b111111111111, 12'b000000000000, 12'b000000000000, 12'b111111110111, 12'b111111111000, 12'b000000001000, 12'b000000000000, 12'b111111110111, 12'b000000000001, 12'b111111111010, 12'b111111111101, 12'b000000001000, 12'b000000000000, 12'b111111110000}, 
{12'b000000101000, 12'b000000010101, 12'b111111110000, 12'b000000000000, 12'b111111101001, 12'b000000000000, 12'b000000001110, 12'b000000000001, 12'b000000001110, 12'b111111111111, 12'b111111110110, 12'b111111111010, 12'b000000001001, 12'b000000000001, 12'b111111111001, 12'b000000001000, 12'b000000100010, 12'b111111110111, 12'b111111101101, 12'b000000000000, 12'b111111111110, 12'b111111110100, 12'b111111111111, 12'b111111111111, 12'b000000000101, 12'b111111101000, 12'b000000000101, 12'b111111111111, 12'b000000000000, 12'b000000000110, 12'b111111111110, 12'b000000000011}, 
{12'b111111111010, 12'b111111110011, 12'b111111111101, 12'b111111110101, 12'b111111111110, 12'b000000000011, 12'b000000000000, 12'b111111111111, 12'b000000000010, 12'b111111111111, 12'b000000000000, 12'b111111110010, 12'b000000000110, 12'b000000000101, 12'b111111111001, 12'b000000011100, 12'b111111111111, 12'b000000000000, 12'b111111111111, 12'b000000000000, 12'b000000010100, 12'b111111100001, 12'b111111111001, 12'b111111111100, 12'b111111111110, 12'b000000001100, 12'b111111111100, 12'b000000000001, 12'b000000011110, 12'b111111011111, 12'b111111101000, 12'b000000000001}, 
{12'b000000000001, 12'b111111111100, 12'b111111111111, 12'b000000000000, 12'b111111010001, 12'b111111011001, 12'b000000000000, 12'b111111111111, 12'b111111101111, 12'b000000000001, 12'b000000000000, 12'b111111111110, 12'b000000000000, 12'b111111111100, 12'b111111111100, 12'b111111111011, 12'b111111110110, 12'b000000010010, 12'b000000000000, 12'b000000000010, 12'b111111111111, 12'b111111111011, 12'b000000000000, 12'b111111111010, 12'b000000001110, 12'b111111011000, 12'b000000001110, 12'b111111111111, 12'b111111111111, 12'b000000001100, 12'b111111111111, 12'b000000001111}, 
{12'b111111111111, 12'b000000000000, 12'b111111111101, 12'b000000000100, 12'b000000000011, 12'b111111101010, 12'b000000000000, 12'b000000000100, 12'b000000100101, 12'b111111111111, 12'b000000000000, 12'b000000000011, 12'b000000010110, 12'b111111111101, 12'b000000000000, 12'b000000000110, 12'b111111111111, 12'b000000000001, 12'b111111111111, 12'b000000000000, 12'b111111101110, 12'b000000000010, 12'b000000000100, 12'b000000000001, 12'b111111111111, 12'b000000001101, 12'b000000000000, 12'b000000001000, 12'b111111100101, 12'b000000000110, 12'b000000011001, 12'b000000000000}, 
{12'b111111101001, 12'b000000001101, 12'b111111101111, 12'b000000000111, 12'b111111111001, 12'b000000000000, 12'b000000011111, 12'b111111110001, 12'b111111101101, 12'b000000001010, 12'b111111110001, 12'b111111111110, 12'b111111111111, 12'b000000010110, 12'b111111111111, 12'b111111101100, 12'b111111111111, 12'b000000011100, 12'b111111100001, 12'b111111111110, 12'b000000010100, 12'b111111101000, 12'b000000000011, 12'b111111111111, 12'b000000010001, 12'b111111011111, 12'b111111101000, 12'b111111110011, 12'b111111111111, 12'b000000000110, 12'b000000000001, 12'b000000001011}, 
{12'b111111111010, 12'b000000000011, 12'b111111111111, 12'b000000001001, 12'b111111111101, 12'b000000001110, 12'b000000000000, 12'b111111111111, 12'b111111111111, 12'b000000000000, 12'b000000000000, 12'b111111111111, 12'b111111111111, 12'b000000100001, 12'b000000000000, 12'b000000001100, 12'b000000000000, 12'b111111110010, 12'b111111111011, 12'b111111111111, 12'b111111111110, 12'b000000000010, 12'b111111111111, 12'b111111110100, 12'b111111111111, 12'b000000010010, 12'b000000010011, 12'b111111111111, 12'b111111111110, 12'b000000000000, 12'b111111111111, 12'b111111111001}, 
{12'b111111111010, 12'b000000000000, 12'b000000010001, 12'b000000000000, 12'b000000000000, 12'b111111111000, 12'b000000000000, 12'b111111001000, 12'b000000001101, 12'b000000000000, 12'b000000000001, 12'b111111101000, 12'b000000000000, 12'b111111110111, 12'b111111111101, 12'b000000000000, 12'b000000000001, 12'b000000000000, 12'b000000000111, 12'b000000000000, 12'b111111111111, 12'b000000010101, 12'b000000011000, 12'b111111110001, 12'b111111110110, 12'b000000001111, 12'b111111101100, 12'b000000000001, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b000000001011}, 
{12'b111111111000, 12'b111111111111, 12'b111111110000, 12'b111111110011, 12'b111111111111, 12'b111111110111, 12'b000000000000, 12'b000000000101, 12'b111111110000, 12'b111111111010, 12'b111111111100, 12'b000000000000, 12'b000000000001, 12'b111111111111, 12'b111111111100, 12'b000000000110, 12'b000000001110, 12'b000000001000, 12'b111111110111, 12'b000000000011, 12'b111111111111, 12'b111111111110, 12'b000000000001, 12'b000000000001, 12'b111111111011, 12'b000000000101, 12'b111111111010, 12'b000000000011, 12'b111111111111, 12'b111111101101, 12'b111111111110, 12'b000000001110}, 
{12'b111111111110, 12'b111111111010, 12'b000000000100, 12'b000000010000, 12'b000000000101, 12'b000000000101, 12'b000000000010, 12'b111111110011, 12'b111111110010, 12'b000000000100, 12'b000000000000, 12'b000000000010, 12'b000000000001, 12'b000000000000, 12'b000000001101, 12'b000000000000, 12'b111111111100, 12'b000000000110, 12'b111111111110, 12'b111111111101, 12'b000000000111, 12'b111111111000, 12'b111111111110, 12'b000000001000, 12'b000000000001, 12'b111111111001, 12'b111111110011, 12'b111111111111, 12'b111111101110, 12'b000000000011, 12'b000000000110, 12'b000000000000}, 
{12'b111111111111, 12'b111111111110, 12'b111111111111, 12'b111111111101, 12'b111111110111, 12'b111111110111, 12'b000000000100, 12'b000000000000, 12'b111111110100, 12'b000000001010, 12'b111111111110, 12'b111111111111, 12'b111111111000, 12'b000000000000, 12'b000000000001, 12'b111111111100, 12'b111111111110, 12'b111111111101, 12'b111111111010, 12'b000000000000, 12'b111111110111, 12'b000000000110, 12'b111111110010, 12'b000000000000, 12'b000000000010, 12'b000000000111, 12'b000000000001, 12'b000000000000, 12'b000000010010, 12'b000000000011, 12'b000000000000, 12'b000000000101}, 
{12'b111111111110, 12'b000000010000, 12'b111111111111, 12'b111111111101, 12'b111111110010, 12'b111111111011, 12'b000000011010, 12'b111111010011, 12'b111111101001, 12'b111111110011, 12'b111111110001, 12'b111111101111, 12'b111111111111, 12'b000000011110, 12'b111111111110, 12'b000000000000, 12'b111111110010, 12'b000000011100, 12'b111111100101, 12'b000000000000, 12'b111111111111, 12'b111111101010, 12'b000000000000, 12'b111111111111, 12'b000000000011, 12'b111111111100, 12'b111111110110, 12'b111111111111, 12'b000000001011, 12'b000000000000, 12'b111111111010, 12'b000000000000}, 
{12'b000000010111, 12'b111111111000, 12'b000000001000, 12'b111111111101, 12'b000000000100, 12'b111111111111, 12'b111111111111, 12'b111111111010, 12'b000000000000, 12'b000000000101, 12'b111111111111, 12'b111111111100, 12'b111111111111, 12'b000000001110, 12'b000000000001, 12'b000000000010, 12'b000000000001, 12'b111111111110, 12'b000000000001, 12'b000000000000, 12'b111111111111, 12'b111111111111, 12'b111111101100, 12'b111111111111, 12'b000000000011, 12'b111111111000, 12'b111111110111, 12'b111111111111, 12'b111111111111, 12'b000000100011, 12'b111111101101, 12'b111111111000}, 
{12'b111111111101, 12'b111111111001, 12'b111111111011, 12'b000000000010, 12'b000000001000, 12'b111111110111, 12'b111111111111, 12'b111111110001, 12'b000000000011, 12'b000000001000, 12'b111111110010, 12'b111111101111, 12'b000000000001, 12'b111111010100, 12'b111111111011, 12'b111111111000, 12'b111111110011, 12'b111111111111, 12'b000000001000, 12'b000000000000, 12'b111111111101, 12'b111111111101, 12'b000000000000, 12'b000000000000, 12'b111111111100, 12'b111111001111, 12'b111111011100, 12'b111111101110, 12'b000000000011, 12'b000000001101, 12'b111111111111, 12'b000000001111}, 
{12'b111111111010, 12'b111111110010, 12'b000000001010, 12'b000000000100, 12'b000000000010, 12'b111111111010, 12'b111111111101, 12'b000000000110, 12'b000000100010, 12'b111111110101, 12'b111111111111, 12'b111111111111, 12'b000000000111, 12'b111111111100, 12'b111111111110, 12'b111111111110, 12'b111111111001, 12'b111111111111, 12'b000000000000, 12'b000000001110, 12'b111111110111, 12'b111111111111, 12'b000000001000, 12'b111111111111, 12'b000000000000, 12'b000000100001, 12'b000000010100, 12'b000000000000, 12'b000000000000, 12'b111111100101, 12'b111111111011, 12'b111111111111}, 
{12'b000000000000, 12'b000000000011, 12'b111111111111, 12'b000000000000, 12'b000000001110, 12'b111111100001, 12'b000000000000, 12'b111111111001, 12'b000000001011, 12'b000000000000, 12'b111111111110, 12'b000000000000, 12'b000000000000, 12'b111111111111, 12'b000000000000, 12'b111111111001, 12'b000000010000, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b000000000000, 12'b111111111111, 12'b000000000000, 12'b111111111111, 12'b000000000000, 12'b111111101011, 12'b000000000011, 12'b000000001011, 12'b111111111111, 12'b000000000110, 12'b111111111111, 12'b000000000100}, 
{12'b111111110011, 12'b000000000000, 12'b111111100001, 12'b000000000000, 12'b111111111100, 12'b111111111101, 12'b111111111111, 12'b111111111010, 12'b111111111101, 12'b111111111011, 12'b000000000011, 12'b000000000001, 12'b111111110100, 12'b000000000000, 12'b111111111111, 12'b111111111111, 12'b000000000100, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111111, 12'b000000010001, 12'b111111111111, 12'b000000000000, 12'b111111111111, 12'b000000010100, 12'b000000001100, 12'b000000000010, 12'b111111111001, 12'b111111111111, 12'b000000000100, 12'b000000000011}, 
{12'b000000000010, 12'b000000000010, 12'b111111111111, 12'b000000000000, 12'b111111100010, 12'b000000000010, 12'b000000000001, 12'b111111111111, 12'b000000000000, 12'b111111110101, 12'b111111111111, 12'b000000000000, 12'b111111110101, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b111111101001, 12'b000000000000, 12'b111111111111, 12'b111111111111, 12'b000000000000, 12'b000000001000, 12'b111111111111, 12'b000000000000, 12'b000000011101, 12'b000000010101, 12'b000000000000, 12'b000000000000, 12'b111111110001, 12'b000000000000, 12'b111111111111}, 
{12'b000000000100, 12'b000000000011, 12'b000000010000, 12'b111111110000, 12'b000000001000, 12'b000000000111, 12'b000000000000, 12'b000000001100, 12'b000000000000, 12'b111111111111, 12'b000000000010, 12'b000000000000, 12'b111111111111, 12'b000000000111, 12'b111111111111, 12'b111111111101, 12'b000000000000, 12'b000000000010, 12'b111111111100, 12'b000000000110, 12'b000000000010, 12'b111111011010, 12'b111111111000, 12'b000000000101, 12'b111111111111, 12'b111111011111, 12'b111111110111, 12'b111111111110, 12'b111111111111, 12'b111111111100, 12'b000000000000, 12'b111111111101}, 
{12'b000000000000, 12'b111111111111, 12'b111111111010, 12'b111111110101, 12'b000000000010, 12'b000000000000, 12'b000000000110, 12'b111111111111, 12'b000000001111, 12'b111111111111, 12'b000000000000, 12'b111111101010, 12'b111111111111, 12'b000000001000, 12'b111111111111, 12'b111111101111, 12'b000000000000, 12'b111111111111, 12'b000000010000, 12'b111111111111, 12'b111111100100, 12'b111111111111, 12'b000000010000, 12'b111111111111, 12'b111111111111, 12'b000000001000, 12'b111111111001, 12'b000000000100, 12'b000000000000, 12'b111111110011, 12'b000000000000, 12'b000000000000}, 
{12'b111111110010, 12'b000000000000, 12'b000000000000, 12'b111111111111, 12'b000000011111, 12'b111111111000, 12'b111111111111, 12'b111111111111, 12'b111111111101, 12'b111111111100, 12'b000000000100, 12'b000000001000, 12'b111111111101, 12'b000000001111, 12'b000000000000, 12'b111111111111, 12'b111111101101, 12'b111111111111, 12'b000000000000, 12'b111111111010, 12'b000000000000, 12'b000000000010, 12'b000000000000, 12'b111111111111, 12'b111111111100, 12'b111111110011, 12'b111111101101, 12'b000000000000, 12'b111111111000, 12'b000000000010, 12'b111111111111, 12'b000000000100}, 
{12'b111111100101, 12'b111111110101, 12'b111111110110, 12'b000000000000, 12'b000000100100, 12'b111111110001, 12'b000000000000, 12'b111111111100, 12'b111111100101, 12'b000000001000, 12'b111111111111, 12'b000000100100, 12'b000000000000, 12'b111111111100, 12'b111111111111, 12'b000000000010, 12'b111111111110, 12'b000000000000, 12'b111111111101, 12'b000000011111, 12'b000000000010, 12'b111111111101, 12'b000000000111, 12'b111111111111, 12'b111111111111, 12'b111111111001, 12'b111111111101, 12'b111111100010, 12'b111111110110, 12'b111111111111, 12'b111111111111, 12'b111111111100}, 
{12'b000000001110, 12'b111111001100, 12'b111111010001, 12'b111111110101, 12'b000000101010, 12'b111111111111, 12'b111111101001, 12'b000000010000, 12'b000000000011, 12'b000000000000, 12'b000000001101, 12'b111111101110, 12'b000000000000, 12'b000000000000, 12'b111111111101, 12'b000000000001, 12'b111111111001, 12'b111111000101, 12'b000000001010, 12'b000000010110, 12'b000000010000, 12'b000000000000, 12'b000000000001, 12'b111111100110, 12'b111111010111, 12'b111111111111, 12'b111111101100, 12'b111111100010, 12'b111111110011, 12'b111111000111, 12'b000000011010, 12'b000000011011}, 
{12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000010000, 12'b111111110100, 12'b000000000001, 12'b000000000100, 12'b111111101001, 12'b000000000010, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b000000001111, 12'b000000000011, 12'b000000000001, 12'b000000000011, 12'b000000010101, 12'b111111110010, 12'b000000000000, 12'b111111110101, 12'b111111111111, 12'b000000010100, 12'b000000000000, 12'b111111111111, 12'b111111011100, 12'b111111111111, 12'b111111110110, 12'b111111111100, 12'b000000000000, 12'b000000001000, 12'b000000000110}, 
{12'b111111111101, 12'b000000001000, 12'b111111101100, 12'b000000000001, 12'b000000001100, 12'b111111111101, 12'b111111111111, 12'b000000001010, 12'b000000000000, 12'b111111111111, 12'b111111111011, 12'b000000000000, 12'b000000000000, 12'b111111111101, 12'b111111111000, 12'b111111111011, 12'b111111111100, 12'b111111111011, 12'b111111111000, 12'b000000000000, 12'b111111111111, 12'b111111111101, 12'b111111111011, 12'b000000011001, 12'b000000000000, 12'b111111101000, 12'b111111111111, 12'b000000000111, 12'b000000000000, 12'b000000000000, 12'b000000010000, 12'b111111111111}, 
{12'b111111111111, 12'b000000000000, 12'b111111111111, 12'b111111110110, 12'b111111001000, 12'b000000000000, 12'b000000000000, 12'b111111111111, 12'b111111011001, 12'b000000000101, 12'b111111111001, 12'b111111111111, 12'b000000000000, 12'b111111101000, 12'b111111111101, 12'b111111111111, 12'b000000000000, 12'b000000000000, 12'b000000000010, 12'b000000010110, 12'b111111111000, 12'b111111101100, 12'b000000000000, 12'b111111101111, 12'b111111111001, 12'b111111110001, 12'b111111111111, 12'b111111111111, 12'b111111111110, 12'b111111100001, 12'b111111111101, 12'b000000001111}, 
{12'b000000000111, 12'b000000001110, 12'b111111111111, 12'b000000001010, 12'b111111110010, 12'b111111111000, 12'b000000000110, 12'b000000000100, 12'b111111111100, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111101011, 12'b111111111111, 12'b000000001001, 12'b111111111000, 12'b000000000010, 12'b111111111111, 12'b111111111111, 12'b000000001101, 12'b111111101011, 12'b000000010001, 12'b000000000011, 12'b000000000000, 12'b000000001101, 12'b000000000000, 12'b111111111101, 12'b111111100111, 12'b111111111000, 12'b111111110101, 12'b000000001011}, 
{12'b000000000000, 12'b000000000000, 12'b111111101000, 12'b111111111111, 12'b000000001101, 12'b111111110110, 12'b111111111111, 12'b111111111111, 12'b000000000001, 12'b000000000000, 12'b000000000000, 12'b111111110010, 12'b000000000110, 12'b000000000000, 12'b000000000000, 12'b000000000010, 12'b111111111111, 12'b111111110110, 12'b000000000001, 12'b000000000000, 12'b111111111101, 12'b111111111110, 12'b000000010010, 12'b111111111111, 12'b000000000000, 12'b111111101101, 12'b111111101011, 12'b000000001111, 12'b111111111111, 12'b111111111111, 12'b000000000001, 12'b000000010010}, 
{12'b111111101010, 12'b111111111111, 12'b111111110010, 12'b000000000000, 12'b111111101001, 12'b000000000000, 12'b111111111111, 12'b111111111011, 12'b111111011101, 12'b111111111110, 12'b000000000000, 12'b111111111111, 12'b111111111111, 12'b000000000000, 12'b111111111111, 12'b111111111100, 12'b111111110110, 12'b111111111001, 12'b000000000100, 12'b111111111111, 12'b111111111110, 12'b000000000000, 12'b000000010101, 12'b111111111111, 12'b000000001001, 12'b000000000101, 12'b111111110111, 12'b000000001101, 12'b111111111101, 12'b000000000000, 12'b111111111111, 12'b000000100101}, 
{12'b111111101011, 12'b000000000001, 12'b000000000011, 12'b111111111110, 12'b000000001111, 12'b111111101100, 12'b111111111111, 12'b000000010000, 12'b000000001010, 12'b000000000000, 12'b111111111111, 12'b111111111011, 12'b111111111010, 12'b111111111011, 12'b111111111100, 12'b000000000101, 12'b111111111111, 12'b000000000000, 12'b000000001001, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000010000, 12'b000000000010, 12'b000000000000, 12'b111111111001, 12'b111111111111, 12'b000000000000, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b000000000100}, 
{12'b111111111111, 12'b000000000000, 12'b111111110010, 12'b111111111011, 12'b000000010010, 12'b111111111111, 12'b111111111011, 12'b000000001111, 12'b111111111100, 12'b000000010010, 12'b000000000101, 12'b111111111000, 12'b000000000000, 12'b000000000000, 12'b111111111111, 12'b000000000001, 12'b111111111011, 12'b111111101111, 12'b000000010001, 12'b000000001001, 12'b000000101000, 12'b000000001100, 12'b000000001111, 12'b111111111111, 12'b000000000000, 12'b000000000000, 12'b000000000011, 12'b000000000101, 12'b111111100101, 12'b111111111111, 12'b111111111111, 12'b111111111111}, 
{12'b000000000000, 12'b111111111010, 12'b111111111001, 12'b000000000000, 12'b111111110000, 12'b000000000000, 12'b000000001100, 12'b000000000110, 12'b000000000011, 12'b111111111001, 12'b000000000000, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111101, 12'b000000001100, 12'b111111111111, 12'b111111111111, 12'b111111101100, 12'b000000000000, 12'b111111110011, 12'b111111111111, 12'b000000000000, 12'b111111111111, 12'b000000000000, 12'b000000000001, 12'b000000000001, 12'b000000001000, 12'b111111111011, 12'b111111111111, 12'b111111100011, 12'b000000000101}, 
{12'b000000011100, 12'b111111111111, 12'b000000000100, 12'b111111111001, 12'b111111111010, 12'b000000000010, 12'b000000001010, 12'b000000000000, 12'b000000100001, 12'b000000000000, 12'b111111111110, 12'b000000000001, 12'b000000000110, 12'b111111111111, 12'b000000000011, 12'b000000000110, 12'b111111111111, 12'b111111100011, 12'b111111111100, 12'b111111111111, 12'b000000000111, 12'b000000000000, 12'b111111111111, 12'b000000000111, 12'b000000000001, 12'b111111101111, 12'b111111111001, 12'b000000001000, 12'b111111111110, 12'b000000010000, 12'b111111111111, 12'b111111110100}, 
{12'b000000000000, 12'b000000000110, 12'b111111111111, 12'b111111111101, 12'b111111101001, 12'b111111111111, 12'b000000000010, 12'b111111111101, 12'b000000001010, 12'b111111111101, 12'b111111111111, 12'b111111111101, 12'b111111111111, 12'b111111111101, 12'b000000000000, 12'b000000010100, 12'b000000000000, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b000000000010, 12'b000000001000, 12'b000000000000, 12'b000000000000, 12'b000000000010, 12'b111111111111, 12'b000000000000, 12'b000000000001, 12'b000000000000, 12'b000000000110}, 
{12'b111111101100, 12'b000000001000, 12'b000000000001, 12'b111111111001, 12'b111111100110, 12'b111111111110, 12'b000000000100, 12'b111111100110, 12'b000000100000, 12'b000000000100, 12'b000000000001, 12'b000000000110, 12'b000000000010, 12'b000000000000, 12'b000000011010, 12'b111111111010, 12'b000000000000, 12'b000000000000, 12'b111111111111, 12'b000000000000, 12'b111111100100, 12'b000000000001, 12'b000000001001, 12'b000000000010, 12'b000000000010, 12'b111111010101, 12'b111111101010, 12'b111111110000, 12'b000000000000, 12'b111111111111, 12'b000000010100, 12'b111111110010}, 
{12'b111111111111, 12'b111111110011, 12'b111111111001, 12'b111111100101, 12'b111111101111, 12'b000000010101, 12'b000000010011, 12'b111111110101, 12'b000000000010, 12'b111111111101, 12'b111111111001, 12'b111111101111, 12'b000000000110, 12'b111111101101, 12'b000000001100, 12'b111111111111, 12'b000000010101, 12'b111111111111, 12'b111111111111, 12'b111111110111, 12'b111111111101, 12'b111111111011, 12'b111111101110, 12'b000000000101, 12'b111111111111, 12'b111111111111, 12'b111111110001, 12'b000000010100, 12'b000000010001, 12'b111111111010, 12'b111111010111, 12'b000000001001}, 
{12'b000000000000, 12'b111111111110, 12'b111111111111, 12'b111111111001, 12'b000000000001, 12'b000000000000, 12'b000000000100, 12'b000000000000, 12'b000000000111, 12'b111111111111, 12'b000000000000, 12'b000000000110, 12'b000000000000, 12'b000000000000, 12'b111111110111, 12'b111111111001, 12'b000000000000, 12'b000000001011, 12'b000000000011, 12'b000000001000, 12'b111111111110, 12'b111111110101, 12'b111111111111, 12'b000000000100, 12'b111111111111, 12'b000000000010, 12'b111111111111, 12'b000000000100, 12'b000000000000, 12'b000000000101, 12'b111111100111, 12'b111111111111}, 
{12'b000000010011, 12'b111111111111, 12'b000000001001, 12'b111111101100, 12'b111111110011, 12'b111111111111, 12'b111111111111, 12'b000000000001, 12'b000000000000, 12'b111111110111, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b111111110111, 12'b000000001001, 12'b111111111111, 12'b111111111110, 12'b000000000000, 12'b000000000111, 12'b111111110011, 12'b000000000111, 12'b000000001000, 12'b000000001000, 12'b111111111111, 12'b000000100011, 12'b111111110110, 12'b000000010111, 12'b111111111100, 12'b111111101000, 12'b111111110100, 12'b000000001000}, 
{12'b111111011101, 12'b111111111110, 12'b111111110110, 12'b111111111111, 12'b000000010000, 12'b111111110100, 12'b111111111100, 12'b000000001111, 12'b000000000110, 12'b111111110000, 12'b000000000000, 12'b111111111110, 12'b111111111111, 12'b000000001000, 12'b111111110000, 12'b111111111111, 12'b000000000000, 12'b111111111111, 12'b111111111110, 12'b000000000000, 12'b111111110011, 12'b111111111111, 12'b000000000000, 12'b111111101010, 12'b000000000100, 12'b000000100111, 12'b000000010110, 12'b111111111101, 12'b111111110101, 12'b111111100011, 12'b000000000000, 12'b111111111100}, 
{12'b000000000001, 12'b000000001101, 12'b000000000001, 12'b111111110110, 12'b000000000000, 12'b111111111110, 12'b000000000000, 12'b000000001101, 12'b000000001101, 12'b111111110111, 12'b000000001000, 12'b000000000001, 12'b111111111111, 12'b111111111111, 12'b111111110101, 12'b000000010000, 12'b111111111101, 12'b111111101011, 12'b000000000111, 12'b111111111111, 12'b111111111111, 12'b000000000111, 12'b111111111011, 12'b111111111111, 12'b111111111100, 12'b000000000101, 12'b111111110111, 12'b000000001000, 12'b111111101000, 12'b000000000101, 12'b111111111111, 12'b000000001010}, 
{12'b111111111101, 12'b000000000000, 12'b000000000101, 12'b000000000000, 12'b111111111100, 12'b111111111111, 12'b000000000110, 12'b111111111111, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000001, 12'b111111111001, 12'b000000000000, 12'b000000000111, 12'b000000000010, 12'b000000000110, 12'b111111111111, 12'b111111111111, 12'b000000001000, 12'b000000001111, 12'b111111111001, 12'b000000000000, 12'b111111111111, 12'b000000000000, 12'b111111100010, 12'b111111111111, 12'b111111111011, 12'b111111111111, 12'b000000100100, 12'b000000000000, 12'b111111110010}, 
{12'b111111111110, 12'b111111111000, 12'b111111111111, 12'b000000000000, 12'b000000000101, 12'b111111111111, 12'b000000000000, 12'b111111111110, 12'b000000000100, 12'b111111111111, 12'b000000000000, 12'b000000000010, 12'b000000010010, 12'b111111111001, 12'b000000000000, 12'b111111001001, 12'b111111111111, 12'b111111111100, 12'b000000000000, 12'b111111111100, 12'b000000000101, 12'b111111110001, 12'b000000000111, 12'b000000000110, 12'b111111111111, 12'b111111010010, 12'b111111110001, 12'b111111111110, 12'b111111111110, 12'b000000011000, 12'b111111111111, 12'b000000001001}, 
{12'b000000000011, 12'b000000000000, 12'b000000001011, 12'b111111111000, 12'b111111111011, 12'b000000001111, 12'b111111110101, 12'b000000000011, 12'b111111101100, 12'b000000000000, 12'b000000000001, 12'b111111111010, 12'b000000000000, 12'b000000000000, 12'b111111110011, 12'b000000011011, 12'b111111110000, 12'b111111111111, 12'b000000000111, 12'b111111111111, 12'b000000000100, 12'b111111100001, 12'b000000010100, 12'b111111111111, 12'b111111111000, 12'b000000011111, 12'b000000001001, 12'b111111110101, 12'b111111110111, 12'b111111011101, 12'b111111111111, 12'b000000000001}, 
{12'b111111111111, 12'b000000000000, 12'b111111111101, 12'b111111101110, 12'b111111111111, 12'b111111100110, 12'b000000000000, 12'b000000010011, 12'b000000001111, 12'b000000000001, 12'b000000000000, 12'b111111111000, 12'b000000010101, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b000000011011, 12'b000000000000, 12'b111111111101, 12'b111111111100, 12'b111111101011, 12'b000000001000, 12'b000000000000, 12'b000000000000, 12'b000000000010, 12'b111111111011, 12'b111111100010, 12'b000000010001, 12'b111111100011, 12'b000000000011, 12'b111111111010, 12'b000000000000}, 
{12'b000000000011, 12'b000000001011, 12'b000000000000, 12'b111111111111, 12'b111111100010, 12'b000000000000, 12'b111111111111, 12'b000000001111, 12'b000000010001, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b111111111111, 12'b000000001010, 12'b111111111001, 12'b111111100100, 12'b111111111101, 12'b111111111001, 12'b111111111001, 12'b111111111011, 12'b111111111111, 12'b111111111011, 12'b111111111110, 12'b111111111111, 12'b000000001001, 12'b111111111111, 12'b000000011101}
};

localparam logic signed [11:0] bias [32] = '{
12'b000001011110,  // 1.474280834197998
12'b000000101100,  // 0.6914801001548767
12'b000001011100,  // 1.4406442642211914
12'b000001011010,  // 1.408045768737793
12'b000000111111,  // 0.9864811301231384
12'b000000110111,  // 0.8636202812194824
12'b111111011000,  // -0.6153604388237
12'b000000011110,  // 0.4839226007461548
12'b000000011111,  // 0.4862793982028961
12'b000000010111,  // 0.37162142992019653
12'b000000011101,  // 0.45989668369293213
12'b000001010011,  // 1.2998151779174805
12'b111110111110,  // -1.016528844833374
12'b111111101001,  // -0.35249894857406616
12'b000000011100,  // 0.44582197070121765
12'b111111111000,  // -0.1119980737566948
12'b111111111011,  // -0.06717441976070404
12'b000000000000,  // 0.00487547367811203
12'b000000001100,  // 0.1946917623281479
12'b111111001110,  // -0.7796769738197327
12'b000000101110,  // 0.7287401556968689
12'b000001101101,  // 1.714877724647522
12'b111110011001,  // -1.5971007347106934
12'b000000000100,  // 0.07393483817577362
12'b000000010100,  // 0.3225609362125397
12'b000000110110,  // 0.8453295230865479
12'b000000111001,  // 0.898597240447998
12'b000000010000,  // 0.2548799514770508
12'b000000111110,  // 0.9735668301582336
12'b000001001000,  // 1.1261906623840332
12'b000000011100,  // 0.44768181443214417
12'b111101101000   // -2.3676068782806396
};
endpackage