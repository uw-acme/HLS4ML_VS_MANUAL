// Width: 8
// NFRAC: 4
package dense_4_8_4;

localparam logic signed [7:0] weights [32][5] = '{ 
{8'b11111111, 8'b00000101, 8'b11111011, 8'b00000001, 8'b11111110}, 
{8'b11110111, 8'b11111111, 8'b00000111, 8'b11111111, 8'b00000000}, 
{8'b00000101, 8'b00000011, 8'b11111111, 8'b11111001, 8'b11111100}, 
{8'b11111001, 8'b11111010, 8'b11111110, 8'b00000100, 8'b00000011}, 
{8'b00000001, 8'b00000010, 8'b00000010, 8'b11111111, 8'b11101111}, 
{8'b00000101, 8'b11111001, 8'b00000010, 8'b11111101, 8'b11111101}, 
{8'b11111001, 8'b00000000, 8'b11111111, 8'b00000010, 8'b00000001}, 
{8'b11111111, 8'b00000100, 8'b11111001, 8'b00000010, 8'b00000010}, 
{8'b00000010, 8'b11111101, 8'b00000000, 8'b11111000, 8'b11111100}, 
{8'b11111111, 8'b11111011, 8'b00000010, 8'b00000110, 8'b00000000}, 
{8'b11111101, 8'b11111101, 8'b00000000, 8'b00001001, 8'b11111011}, 
{8'b00000010, 8'b00000011, 8'b11111010, 8'b11111111, 8'b00000001}, 
{8'b00000000, 8'b00000010, 8'b00000000, 8'b11111100, 8'b11110110}, 
{8'b00000010, 8'b00000001, 8'b00000110, 8'b11111110, 8'b11111001}, 
{8'b00000001, 8'b11111111, 8'b11111010, 8'b11111111, 8'b00001000}, 
{8'b11111000, 8'b11111100, 8'b11111100, 8'b00000110, 8'b00000000}, 
{8'b00000101, 8'b11111101, 8'b11111101, 8'b11111100, 8'b11111111}, 
{8'b00000011, 8'b11111111, 8'b11111001, 8'b11111111, 8'b00000001}, 
{8'b00000100, 8'b00000000, 8'b11111100, 8'b00000000, 8'b11111001}, 
{8'b00000011, 8'b11111110, 8'b11111100, 8'b00000011, 8'b00000001}, 
{8'b00000001, 8'b11111111, 8'b00000100, 8'b11111001, 8'b11111111}, 
{8'b00000000, 8'b00000001, 8'b00000111, 8'b11110111, 8'b11110110}, 
{8'b11111110, 8'b00000001, 8'b00000010, 8'b11111010, 8'b00001000}, 
{8'b11111111, 8'b00000010, 8'b00000100, 8'b00000000, 8'b11110110}, 
{8'b11111101, 8'b00000101, 8'b11111100, 8'b00000000, 8'b00000110}, 
{8'b00000000, 8'b00000100, 8'b00000000, 8'b11110100, 8'b00001000}, 
{8'b11111000, 8'b11111100, 8'b00000011, 8'b00000011, 8'b00000011}, 
{8'b00000000, 8'b00000011, 8'b11111111, 8'b11111101, 8'b00000000}, 
{8'b11111110, 8'b00000011, 8'b11110111, 8'b00000010, 8'b11111101}, 
{8'b11111111, 8'b00000010, 8'b11111101, 8'b11111001, 8'b00001001}, 
{8'b00000111, 8'b00000001, 8'b00000101, 8'b11110110, 8'b11111010}, 
{8'b11111111, 8'b11111001, 8'b00000101, 8'b00000001, 8'b00000010}
};

localparam logic signed [7:0] bias [5] = '{
8'b11111111,  // -0.06223141402006149
8'b11111110,  // -0.06270556896924973
8'b11111110,  // -0.07014333456754684
8'b00000001,  // 0.0820775106549263
8'b00000011   // 0.2155742198228836
};
endpackage