//Width: 37
//Int: 13
package dense_3_gen;

localparam logic signed [36:0] weights [32][32] = '{
{37'b1111111111111111100110110110011011011, 37'b1111111111111100100000001001001111111, 37'b1111111111111100110000010011010001101, 37'b1111111111111110011110011111100111100, 37'b0000000000000010101111101101010101000, 37'b0000000000000000010110011110010110111, 37'b1111111111111111111001011100011010010, 37'b1111111111111111111111100101101110001, 37'b1111111111111111111111111111000001011, 37'b1111111111111111111111111010001001111, 37'b0000000000000001000000100011011101010, 37'b1111111111111011110010001111101010001, 37'b1111111111111111100001011100001110010, 37'b0000000000000110110001101101011111110, 37'b1111111111111110000100010110010110011, 37'b1111111111111000100010011101010010001, 37'b1111111111111111101101011000100100000, 37'b0000000000000000111001000011101000110, 37'b0000000000000011011110101100110101011, 37'b1111111111111101001101101011010001101, 37'b1111111111110111011110011000010001000, 37'b1111111111111111101000011111011010110, 37'b0000000000000000011001001101011000111, 37'b1111111111111100110001100000111011011, 37'b0000000000000000000000000110011110110, 37'b0000000000001000000110011110000100110, 37'b1111111111110100010110010010110111100, 37'b1111111111111110001110100000111101101, 37'b1111111111111100111001000101000011011, 37'b1111111111111110110011001010000111001, 37'b0000000000000011011000100111000111110, 37'b1111111111111110101110011010101001001},
{37'b0000000000000101111110110100001100011, 37'b0000000000001101110101110001010011110, 37'b0000000000000011001101110111000111110, 37'b1111111111111010101111010001001010011, 37'b0000000000000001111101000101011100000, 37'b1111111111111101110100000010011010111, 37'b1111111111111111001000011101110111000, 37'b0000000000001000101110000001011001110, 37'b0000000000000000000011000011111000000, 37'b1111111111111111111111111100100111101, 37'b1111111111111111101111101111110000100, 37'b1111111111111011010010110101110011000, 37'b1111111111111110011000111001010001000, 37'b0000000000000100010100101011011101111, 37'b1111111111101111001001110101111010100, 37'b1111111111111100001110101110000001100, 37'b1111111111111111111111111110011100111, 37'b1111111111111111111011110000101010010, 37'b1111111111111111100101000010110011100, 37'b1111111111111110101011111000010110100, 37'b1111111111111101111011101101100100000, 37'b1111111111111101110011000001011010001, 37'b0000000000000000001000110101101011111, 37'b1111111111111111111111001010101100010, 37'b1111111111111111111100101101101011001, 37'b1111111111110111011011000100110011000, 37'b0000000000000000000110000000011110010, 37'b0000000000000011110001001000100110011, 37'b1111111111111111011111100110100000100, 37'b1111111111111010011110110101011010001, 37'b0000000000000000000001011000101001110, 37'b0000000000000000010011011000010111011},
{37'b1111111111111000000111100100011101100, 37'b0000000000000001011110010011111111100, 37'b0000000000000000000101011111101111011, 37'b0000000000000010100101001110000011000, 37'b1111111111111010111101010001011111010, 37'b0000000000000000000000010000101001101, 37'b0000000000000000000000110110001100110, 37'b1111111111111001010010010111001010111, 37'b0000000000000100010010011000111001011, 37'b1111111111111101111001110111000101110, 37'b1111111111111101111011001010100000001, 37'b1111111111110100000110101101110010100, 37'b1111111111111101100000110011100110111, 37'b0000000000000100000101100110000010010, 37'b0000000000000010000111000101001010100, 37'b1111111111111111111111001001000010001, 37'b1111111111111111000101011100110100101, 37'b1111111111111111110011111001011010011, 37'b1111111111111001011110111101101111010, 37'b0000000000000000000001100110011000001, 37'b0000000000000000111111110100111000101, 37'b0000000000000000100011010100101101110, 37'b0000000000000001101011000111000010000, 37'b0000000000000111000010100110101000100, 37'b0000000000000000010011011000001111101, 37'b1111111111111001101100011110110111100, 37'b0000000000000110001000111000010001100, 37'b0000000000000000000000010110101110000, 37'b0000000000000001010100111010011110001, 37'b1111111111111111110100101111001111001, 37'b0000000000000000000000011111001000011, 37'b0000000000010010001001101010100101100},
{37'b0000000000000110101100111001101001010, 37'b1111111111111111111111111110010000000, 37'b1111111111111110011100011111011100000, 37'b0000000000001010011110000011100011110, 37'b0000000000001001110100110001110101010, 37'b0000000000000000000000001010111011111, 37'b0000000000000000100101101110100010110, 37'b0000000000000110100000101011011100111, 37'b1111111111111100110101010011100100111, 37'b1111111111111111111111111010000111010, 37'b1111111111111001011010011111101101011, 37'b0000000000000000111101010001011000100, 37'b0000000000000010001000011101100001110, 37'b1111111111111010000001010100010011100, 37'b0000000000000000101111111001000110110, 37'b1111111111111110101110001011100101110, 37'b1111111111111111111111111011110010110, 37'b1111111111111101000101100110111011101, 37'b0000000000000000010011101100010111001, 37'b0000000000000000011100010000101001000, 37'b0000000000000000001000001000100011100, 37'b1111111111111111011010101001000101001, 37'b0000000000001001100011001010110001010, 37'b0000000000000101011111000110111011000, 37'b0000000000000101010001010000001011111, 37'b0000000000000011111110001001001011100, 37'b0000000000000101011101110010101111100, 37'b0000000000000000000000001110010111010, 37'b1111111111111111000011100101011101010, 37'b0000000000000111001111111100111110111, 37'b0000000000000011111111100010100011000, 37'b1111111111111110100110000110011101111},
{37'b0000000000001000000000010000000000000, 37'b1111111111111111010000001011001001010, 37'b1111111111111010011101000111001101110, 37'b1111111111110011111110011011110101000, 37'b0000000000000111101000111010001100100, 37'b0000000000000000000000001000010100100, 37'b1111111111111001011011111111111111000, 37'b1111111111111011011110100110101001001, 37'b1111111111111111010000010100011001001, 37'b1111111111110011000011010111111110010, 37'b1111111111101110010100101010111011100, 37'b0000000000000111100100000011001001110, 37'b0000000000001010101100110100111101110, 37'b0000000000001000010111111001000101100, 37'b1111111111110110110011001011000110100, 37'b1111111111110011100110011010000001010, 37'b0000000000000000000000000100000110101, 37'b1111111111111101101111001100100011111, 37'b0000000000000011001101100010111101100, 37'b0000000000000010001110000010101001000, 37'b1111111111111100111111000110111000000, 37'b1111111111111111111001011111011110001, 37'b0000000000001011100010111111110100010, 37'b1111111111101010000000010001001001100, 37'b0000000000000001011010001000101111111, 37'b1111111111110101011101101000001110010, 37'b0000000000000001000011000110110101100, 37'b1111111111111100000001111010011011111, 37'b1111111111111011001110011001111010100, 37'b1111111111111111111111101011011010011, 37'b0000000000000001000111101010111101000, 37'b0000000000001001010010011101110111100},
{37'b0000000000000000101100001110101110100, 37'b1111111111111111010101101010110010111, 37'b1111111111111011000101100110111011011, 37'b1111111111111011110101011101011101010, 37'b0000000000000101111100101001000010111, 37'b0000000000000000000000001010111110110, 37'b1111111111111011100001100001101000011, 37'b1111111111111101110100100111100001111, 37'b1111111111111001001001100100101101101, 37'b1111111111111110111110011010000110001, 37'b1111111111111111111111100001110010100, 37'b0000000000000010100100001010100001100, 37'b0000000000000000000000000000110110100, 37'b0000000000000101101110010111011001010, 37'b1111111111110111111010000101101001100, 37'b1111111111111101111101010010101010101, 37'b0000000000000001011011001100001100010, 37'b1111111111111011010011111110100001011, 37'b1111111111111100110101101110110010001, 37'b1111111111111111111111111011100001001, 37'b0000000000000000001100011110011110110, 37'b0000000000000100110010110111111000111, 37'b0000000000000111011110001111001010010, 37'b1111111111111111110101000100001111011, 37'b1111111111111111111111100100001100110, 37'b0000000000000110011010010101100111101, 37'b1111111111110111001101010011111100100, 37'b1111111111111111111111111000010011000, 37'b1111111111111100001101110011101100001, 37'b1111111111111111011010010010010110111, 37'b1111111111111111111100110000100100010, 37'b0000000000000000000110101000100000100},
{37'b0000000000000001000010101000010100110, 37'b1111111111111010101011100111100100110, 37'b0000000000000001101110111101111100101, 37'b1111111111111111011000100110111100110, 37'b1111111111111111111000010010101100100, 37'b0000000000000010011011000011001010010, 37'b1111111111111110010011011111011000011, 37'b1111111111110101001010101011000111010, 37'b1111111111111111111111111010001110110, 37'b1111111111111100101010101001111010010, 37'b1111111111111000101100010011100001101, 37'b0000000000000111100011100011110101101, 37'b0000000000000000000111010011110000110, 37'b0000000000001010111100110011101000100, 37'b0000000000001101010000100101000101110, 37'b0000000000000000000010101010101001110, 37'b1111111111111111111111111111001111111, 37'b1111111111111010111101001000001101111, 37'b1111111111111111000000100101101111111, 37'b0000000000000100010111111011011010000, 37'b1111111111110011111111111011111010100, 37'b0000000000000010011111101110010101010, 37'b0000000000000101001110001000011001000, 37'b0000000000000000010011011110000010100, 37'b0000000000000010011001101111010100100, 37'b0000000000010011111001001000100100000, 37'b1111111111111001101100011011010011111, 37'b1111111111111110100011001100101010000, 37'b1111111111111100111101100100000111101, 37'b0000000000000111110010110001010011101, 37'b1111111111111111001101101000100001011, 37'b1111111111111101010010100100000010111},
{37'b1111111111110110011101011011010110100, 37'b0000000000000000011000011000100110000, 37'b1111111111110101111011101111000000110, 37'b0000000000000110111101101001011010101, 37'b0000000000010000011100101000010000100, 37'b0000000000000001110110111000111011111, 37'b0000000000000000000011111010110110001, 37'b0000000000000000110000010100101100100, 37'b1111111111111111111111111110000010100, 37'b0000000000000010000011000011100101110, 37'b0000000000010100110100010010011001000, 37'b1111111111111111111111101101111011000, 37'b0000000000000110000110010111101110110, 37'b0000000000001001111101111001001001110, 37'b0000000000001100010011000010101000000, 37'b0000000000010000110011010100001100000, 37'b0000000000000000000000000011000001101, 37'b1111111111111000010110011001110110101, 37'b0000000000000101011000010110010000001, 37'b1111111111111111111010011000001110101, 37'b1111111111110101110010110110000100100, 37'b1111111111111100010111101100111011100, 37'b0000000000000000001101110011000011100, 37'b1111111111111110101011001110000000011, 37'b1111111111110111111110101000000110100, 37'b0000000000011110000000100011111101100, 37'b1111111111111100011111001000001011000, 37'b0000000000000000000000000011101010000, 37'b0000000000000000000000000011000000010, 37'b0000000000001110001000001110111110010, 37'b0000000000000001011010110010110010111, 37'b0000000000000110010001001011111101000},
{37'b0000000000000110110000011010001111110, 37'b1111111111111111101100000111000011001, 37'b0000000000000000000000010010010000101, 37'b1111111111111111010011101000011011111, 37'b0000000000000001010011100011101101010, 37'b1111111111111111011001000001001001010, 37'b1111111111111111111111101110010011000, 37'b0000000000000010100000101010110010101, 37'b0000000000000011011000011100000011000, 37'b1111111111111011100111011100011111100, 37'b0000000000000010001111011010011010110, 37'b0000000000000010111111111000111100110, 37'b0000000000000000001100001001000100101, 37'b0000000000000101010100110000111101111, 37'b1111111111111100011001100010111110101, 37'b1111111111110011001111111011111000110, 37'b0000000000000000000000000011001011110, 37'b1111111111111111110001101101101101100, 37'b1111111111111111100100101011011101101, 37'b1111111111111000000001011110000000000, 37'b1111111111111111111110110111010111101, 37'b0000000000000000000000000110000100110, 37'b1111111111111100110000011001011100100, 37'b1111111111111111110001100010000100000, 37'b1111111111111110011110101111101110000, 37'b0000000000000010011111100000010000111, 37'b0000000000000101111110101011000011111, 37'b1111111111111110000101101001111000100, 37'b1111111111111111001101101101110100110, 37'b1111111111111111010110110010110010010, 37'b0000000000000000011011101011100110111, 37'b1111111111111001101110001011011000100},
{37'b1111111111111101001010000101000110111, 37'b0000000000000110001001101001001010101, 37'b0000000000000000000000000111100011110, 37'b0000000000000000000000000010111101111, 37'b0000000000001100101011010100001010100, 37'b0000000000000101001001111101110100100, 37'b1111111111111111111111111110011001010, 37'b1111111111110111000111100111100101010, 37'b0000000000000001111000101100110001010, 37'b1111111111110100110101101011010010000, 37'b1111111111101001100011001110110111100, 37'b1111111111111111111111111011100111100, 37'b0000000000000000000000010101001101001, 37'b0000000000000110110111010000011110100, 37'b0000000000000001110001101000111111110, 37'b0000000000000000000000000101111011000, 37'b1111111111111010101111101001111001111, 37'b0000000000000000000000010111011111010, 37'b0000000000000000000110111001001100100, 37'b0000000000000000111110000100100011110, 37'b0000000000000011111001101010001110010, 37'b1111111111111111100101111100011000011, 37'b1111111111111010001111001011110111011, 37'b0000000000000000001000011011100011100, 37'b1111111111111111110100011011000000100, 37'b0000000000010001010011011000010110100, 37'b0000000000000101001110011101101110100, 37'b1111111111111111111111100111010011010, 37'b1111111111111110110111011101001010101, 37'b0000000000001010101100010110100000000, 37'b1111111111111111010111001110100000100, 37'b1111111111111110100110010111001110000},
{37'b1111111111110111101000011110110101010, 37'b0000000000000010110011011111101100101, 37'b1111111111111111011100011111101011111, 37'b1111111111111111111111111010110011010, 37'b1111111111111100000011111001111010110, 37'b1111111111111001111101010010001010011, 37'b0000000000000000110001001101010101010, 37'b0000000000000010010011101011100010010, 37'b1111111111111111111111111110111000100, 37'b1111111111111101010000101110101100110, 37'b1111111111110110110101101010111010100, 37'b0000000000000011001101101001000101000, 37'b0000000000000100110111011100111000001, 37'b0000000000000000000000000010001011010, 37'b0000000000001101011011000110100010010, 37'b1111111111110111000000110001111001000, 37'b0000000000000001101010011101000110110, 37'b1111111111111001101111100110000101001, 37'b0000000000000100100000110000100111011, 37'b1111111111111111111111110001111010001, 37'b1111111111111111011000100011110111100, 37'b0000000000000001000111111101101111100, 37'b0000000000000001111101101000001100011, 37'b0000000000000000000000001000001000001, 37'b1111111111111000000110011100110111001, 37'b0000000000000000011111110111110111110, 37'b1111111111110111000011110010110110010, 37'b1111111111111111010111010011000100000, 37'b1111111111111111111111110001111110100, 37'b0000000000001010110011111110010110000, 37'b1111111111111100111101010111101110001, 37'b0000000000000000000000010010001101100},
{37'b1111111111111111111111111011110010011, 37'b0000000000000001110101100110101001001, 37'b0000000000000000000000010001110010000, 37'b0000000000000110010000101011010010000, 37'b1111111111111110001000000110010100011, 37'b1111111111111111010011111000010111100, 37'b0000000000000000111011111100111011100, 37'b1111111111111111111010000010011010000, 37'b1111111111111111010000100111001100000, 37'b0000000000001010010000000001111110110, 37'b0000000000001011001011111000011101000, 37'b0000000000000000000000101100100110010, 37'b1111111111111010101011011111001101110, 37'b1111111111110100110000111000101001000, 37'b1111111111111111001100000101100011100, 37'b0000000000000000000000001010001001100, 37'b0000000000000000000000001010000100010, 37'b1111111111111110111110110001000101111, 37'b1111111111111000011000000101010010001, 37'b0000000000000110000111100010001100100, 37'b0000000000000000000010001001111001110, 37'b0000000000000101111011111001000101011, 37'b1111111111111111111111110000001100101, 37'b0000000000001000111111111101111100110, 37'b0000000000000001111110101101110010101, 37'b0000000000000100111001101100001011001, 37'b0000000000000111010010011110111010110, 37'b1111111111111111001011000010101100111, 37'b1111111111111001101111001011101101001, 37'b1111111111111000111100110010000101001, 37'b1111111111111111111010110100010110011, 37'b1111111111110101010011000010111100110},
{37'b1111111111111100011000001111111001101, 37'b1111111111111111111111111100000010110, 37'b0000000000000001111010001001100000101, 37'b1111111111111001010011000000011001011, 37'b0000000000000001011000001100101100101, 37'b1111111111111111111111111001001010111, 37'b1111111111111100100001100111100011001, 37'b1111111111111111110110001001111000100, 37'b1111111111111101111111100110001011101, 37'b0000000000000000100110000011100011100, 37'b0000000000000001001111110101110110100, 37'b1111111111111110110110110111010100101, 37'b0000000000000000010000111001010000101, 37'b0000000000000011000000001001010101000, 37'b1111111111110101111111111101100011100, 37'b1111111111111100000101011110000101101, 37'b0000000000000011101001101001001101101, 37'b1111111111111101001010110111010110010, 37'b0000000000000000000000000101001010100, 37'b1111111111111111100110010010101110101, 37'b0000000000000011000101100111110011010, 37'b0000000000000000001000001101000101001, 37'b1111111111111111100000001001100100010, 37'b0000000000000000101011100000111010111, 37'b0000000000000100010011111011111100001, 37'b1111111111111110010101100110101100111, 37'b0000000000000000000000001100000010101, 37'b1111111111111000110001011100111100101, 37'b1111111111111100110111100100100001101, 37'b1111111111111111111000110101001111111, 37'b0000000000000010110001100011000000010, 37'b0000000000000000000000010111011111011},
{37'b1111111111110111101011110000100110110, 37'b0000000000000110101110011101110001000, 37'b1111111111111111111111111100011111000, 37'b1111111111111111111001001011110010111, 37'b1111111111111111110110001000001000001, 37'b0000000000000010110011100010101101011, 37'b1111111111111111111111110000010111010, 37'b0000000000001100010110100111000101100, 37'b1111111111111111110000110111111110111, 37'b1111111111111111111111111101011110000, 37'b0000000000000011010010110000010001100, 37'b0000000000000000101001111110010100000, 37'b0000000000000000000110101010011100000, 37'b0000000000000000000000001110110111101, 37'b0000000000000001111100101100100111100, 37'b0000000000000101010010000110110111000, 37'b0000000000000010110110011100001100110, 37'b0000000000000010101010101110010011001, 37'b1111111111111111110111010001110110001, 37'b0000000000000100111010100111111100001, 37'b0000000000000001100111000100000110111, 37'b0000000000000000101001011111010001011, 37'b1111111111111111110111001100000001001, 37'b0000000000000100000100000101000010010, 37'b1111111111111110011010000000111101101, 37'b1111111111111010100100111110100101101, 37'b1111111111111110100001011011011010100, 37'b1111111111111111111111111100011011111, 37'b0000000000000001101000000010110011010, 37'b0000000000000000011110011010100000100, 37'b0000000000000011001000000100000111100, 37'b0000000000000111101010101001001000010},
{37'b1111111111111111101100111000000001111, 37'b1111111111111001110001010111010110100, 37'b0000000000000000110100111000011011010, 37'b1111111111111111111111000000010110000, 37'b0000000000001110101010000101010101100, 37'b1111111111111100101011101010111011001, 37'b1111111111110110110110101101010100010, 37'b0000000000000000000000001101000011000, 37'b0000000000000000000000000111110100000, 37'b1111111111111111100101100101010011011, 37'b0000000000000000110001100111011110100, 37'b0000000000000110111111001111000011011, 37'b0000000000000101001001101011101000100, 37'b0000000000000000001010111011101011000, 37'b0000000000000000100010001001010001101, 37'b1111111111111101001101000100110110111, 37'b0000000000000000100010001001011110110, 37'b1111111111111111011001001000101010011, 37'b0000000000000000000000000110100101100, 37'b0000000000000001001101001100000011011, 37'b1111111111111111011001101010101111010, 37'b0000000000000000010011100111110011110, 37'b0000000000000100010000101001100111000, 37'b0000000000000000100101110001110110100, 37'b1111111111111111110011101010000110111, 37'b1111111111111001011001011000001101110, 37'b0000000000000011010000000101010111000, 37'b1111111111111111111111111011111111011, 37'b1111111111111111111111101001100011001, 37'b1111111111111110010011001001000101001, 37'b1111111111111111101010000010001100011, 37'b1111111111111110111111111011010100111},
{37'b0000000000000000000111010001101110100, 37'b1111111111111110111111001100011101001, 37'b1111111111111101111110111000111011101, 37'b1111111111111100100000000000110110101, 37'b1111111111110111010000010011001101110, 37'b0000000000001001110000000100101010000, 37'b0000000000000000000000001111010010000, 37'b0000000000000010101100111110110100000, 37'b0000000000000100100101111000001100100, 37'b0000000000000000001101001000101100010, 37'b1111111111111111011101010111000000001, 37'b0000000000000111100111000110000101101, 37'b0000000000000011100101001110100100101, 37'b1111111111111010001001101010010010101, 37'b1111111111111101011001110000000011100, 37'b1111111111111111010101110110101000011, 37'b1111111111111001101000000000100010111, 37'b1111111111111111101110001110010100100, 37'b0000000000000000000000001101100011111, 37'b1111111111111111111011010100011101111, 37'b0000000000000010011111101110100010010, 37'b1111111111111101110011111110011101000, 37'b0000000000000000000000000010110010100, 37'b0000000000000001001110110100100010000, 37'b1111111111111111111111111010100010001, 37'b1111111111111010100010000110100101001, 37'b0000000000000010100000011110101001000, 37'b0000000000000000000000011010010101011, 37'b0000000000000000101101101111111101110, 37'b0000000000000000001011001110011101011, 37'b1111111111111010111100010110011101110, 37'b0000000000000000010101010001101111111},
{37'b1111111111111100110111001110010010110, 37'b1111111111111101011110110110111100011, 37'b0000000000000001001110010001001101100, 37'b1111111111111110000000111010100011001, 37'b1111111111111110100100000001100110001, 37'b0000000000000001110110111110100111110, 37'b1111111111111111111010110000011000000, 37'b0000000000000000100011110001011000000, 37'b0000000000000010000110001000101111010, 37'b1111111111111111111111101000101110110, 37'b0000000000000001111110101110001000110, 37'b1111111111111101111101101010000011001, 37'b1111111111111111110110000100001110011, 37'b1111111111111111111111110100001000100, 37'b0000000000000001101001111010011111011, 37'b1111111111111111111111111010011000010, 37'b0000000000000111110100001110001101011, 37'b1111111111111111101110001111010111010, 37'b0000000000000011111110000000000010100, 37'b1111111111111101010010001010111000110, 37'b0000000000000010100010000011001110110, 37'b0000000000000001000000010110000001001, 37'b0000000000000001010110011010100100110, 37'b0000000000000000100101001001011001010, 37'b1111111111111110101100101000110100100, 37'b1111111111111011100010100001011110110, 37'b1111111111111011110110101101110111110, 37'b0000000000000001101110100000000110010, 37'b1111111111111110101010010010110000011, 37'b0000000000000000000000100101100010100, 37'b1111111111111111100011111101001001011, 37'b0000000000000011101101101010010110010},
{37'b1111111111111111111111111010001011001, 37'b1111111111111001100001011100111011110, 37'b1111111111111001101001111100100010101, 37'b1111111111111111111111111001101110001, 37'b0000000000001010000110011111111101010, 37'b1111111111111110100011000100000101011, 37'b0000000000000000000000001010011010010, 37'b0000000000000111101110111001010100110, 37'b1111111111111101101000111110010100001, 37'b0000000000000000000000000100101110001, 37'b1111111111111001010100010001010101011, 37'b1111111111111000001010000101110100000, 37'b0000000000000111001011000010111111111, 37'b0000000000000010011010110001101000000, 37'b1111111111111110000011110010000000000, 37'b1111111111111011100111101101011100110, 37'b0000000000000010110000100010100110111, 37'b0000000000000000000000011101100010010, 37'b1111111111111100001100100100100101111, 37'b0000000000000000011011001100110001110, 37'b0000000000000001000111001100101010011, 37'b1111111111111110100101011110101101111, 37'b0000000000000100100010110101100110000, 37'b1111111111110000010100110010111010000, 37'b0000000000000000101001111110110011100, 37'b0000000000000011110100110010110100111, 37'b1111111111111111010101110111011101010, 37'b0000000000000000001111010001001001111, 37'b1111111111111100010001001000110100101, 37'b1111111111111111111111110110110000000, 37'b1111111111111100110010000000100000011, 37'b1111111111111111100111010101100111111},
{37'b0000000000000011011001101101110000010, 37'b0000000000000101100001011101110001011, 37'b0000000000001000110011111111010100000, 37'b1111111111111100101110100101100010011, 37'b0000000000000110101010000101101000110, 37'b0000000000000100111001101011110100111, 37'b0000000000000000000000100000101101010, 37'b0000000000000111010010011000010110110, 37'b0000000000000101101101101111101110100, 37'b1111111111111110010010100111000000111, 37'b0000000000001011001110011110100000000, 37'b1111111111111010011010011010011001010, 37'b0000000000001001111100010000110011000, 37'b0000000000000111001001000110001111010, 37'b1111111111101110110101010001101100000, 37'b1111111111111111111111000000101001100, 37'b0000000000000000000000000100001000111, 37'b0000000000000000000101111001100001000, 37'b0000000000000100001010001010011011101, 37'b1111111111110111111100101111000101110, 37'b0000000000000011100010111111010100110, 37'b1111111111111100100110111111110001011, 37'b1111111111111000001001111110000011110, 37'b1111111111111101011111011000100011001, 37'b0000000000000101010001010001100010101, 37'b1111111111110101011100011001101011010, 37'b1111111111111010101110010101001010000, 37'b1111111111111111010101110100100001101, 37'b1111111111111111111111110110000011110, 37'b1111111111110110111110001011001000110, 37'b0000000000000110010100111110011101111, 37'b0000000000000000000000011001000101100},
{37'b1111111111111111001101100001011101000, 37'b0000000000000000000000101111001011011, 37'b1111111111111111111111111100110000010, 37'b1111111111111111111111111110101100100, 37'b1111111111111010011000011010010001010, 37'b0000000000000000001001011010100101011, 37'b0000000000000000001000011100010000010, 37'b1111111111111111110000100111111100110, 37'b1111111111111111100111001111100110001, 37'b1111111111111111010000111011111111001, 37'b0000000000000010001110010100100101001, 37'b1111111111111111111111001111110011111, 37'b0000000000000001010100111010101111100, 37'b1111111111111010100001100111001101111, 37'b0000000000000001101101011111010001111, 37'b1111111111111111111111010001010000010, 37'b0000000000000010010000000110011010100, 37'b0000000000000111001010011011010011101, 37'b1111111111111010010110110101010011101, 37'b0000000000000000110101001000110001000, 37'b1111111111111110011010100011110011001, 37'b0000000000000010000011101110010010100, 37'b0000000000000011000010101100000101100, 37'b1111111111111110101000101100100010111, 37'b1111111111111011111110110001000111010, 37'b0000000000000000010101000101100001001, 37'b0000000000001101010001001101011010000, 37'b1111111111111111100111001101110011100, 37'b1111111111111111110000010110011100010, 37'b0000000000000101001100000110011011001, 37'b0000000000000000000000001101010110000, 37'b0000000000001101110010101101111101010},
{37'b1111111111110111101001111001100010010, 37'b0000000000000000100101000001010000011, 37'b1111111111111100100010011111001010101, 37'b0000000000000110001000000111111100010, 37'b0000000000000001110000010110100100011, 37'b1111111111111111011111101000010111011, 37'b1111111111111111111111111101111001110, 37'b1111111111111111111111111111010011000, 37'b1111111111111011001001100111011110000, 37'b1111111111111111011110001111001110111, 37'b0000000000000000000000001001010110011, 37'b1111111111110111000111011001010100000, 37'b0000000000000000001100110101101110010, 37'b1111111111111111010111010010010101001, 37'b1111111111111111111101011111111010001, 37'b1111111111111111111111110011110110001, 37'b1111111111111110001000100010101001111, 37'b0000000000000000000101100100100011111, 37'b0000000000000000000011001110111101010, 37'b0000000000000010100010011111111111011, 37'b0000000000000000010001111100100000010, 37'b0000000000000000000000000010000110010, 37'b0000000000000000000000001000110011111, 37'b1111111111111111110111101101111001111, 37'b0000000000000000000000010011000001101, 37'b0000000000000000010010110000001111001, 37'b0000000000001001010011010011111001000, 37'b1111111111111111111111111101111000100, 37'b1111111111111111111111110100101111111, 37'b1111111111111111010110010010100111001, 37'b0000000000000010110011010001000111011, 37'b1111111111111111100101111010010011011},
{37'b1111111111111111111110011000011000000, 37'b1111111111111101100101000000011000001, 37'b0000000000000011010001001101001001000, 37'b0000000000000000101000111011001010011, 37'b1111111111111010000011010110110111110, 37'b0000000000000000000000100111110011111, 37'b0000000000000100100100110100000101011, 37'b1111111111111111111111110110100100011, 37'b0000000000000000000000000011011100000, 37'b1111111111111110011011000010101000101, 37'b0000000000000001110101101111010001000, 37'b0000000000000000010011011101101010111, 37'b0000000000000101001011010101101010000, 37'b1111111111110111001110100111001100010, 37'b1111111111111110011111001110100000001, 37'b1111111111111111101110011001001000111, 37'b0000000000000011011101010111000001110, 37'b1111111111111001110110101110011110101, 37'b0000000000000000010101110000000100001, 37'b1111111111110011111011010000110001110, 37'b1111111111111111101100101010101110110, 37'b1111111111111110000110001101111001001, 37'b1111111111111111010110101110000100000, 37'b0000000000000100101110110001110010011, 37'b1111111111111110110011101110000110110, 37'b1111111111111011100000001110010111110, 37'b0000000000000001011100100001100111100, 37'b0000000000000000000000010100010110110, 37'b0000000000000110010101010100111101100, 37'b0000000000001000010111110011111001000, 37'b1111111111111010110000000100001010000, 37'b1111111111111000110100000000011110001},
{37'b0000000000000001000101000100101101000, 37'b0000000000000000011010001001011101100, 37'b1111111111111001010111111110001000000, 37'b1111111111111111000101111000001110100, 37'b1111111111111111111111111001000100010, 37'b0000000000000000000010001110110010111, 37'b0000000000000001101100110100001000100, 37'b0000000000000110100101001111001011100, 37'b0000000000000000000000000101000011111, 37'b0000000000000000010100110001110110010, 37'b0000000000000001000111101101011001000, 37'b1111111111110111010111101011000000110, 37'b1111111111111110111011110100010000111, 37'b1111111111110110010101110001001011100, 37'b0000000000000111101100011000000111001, 37'b0000000000000000000000011010101000100, 37'b1111111111111111111111001101101110001, 37'b1111111111110101101111110101111100000, 37'b1111111111111111111111101111001000011, 37'b1111111111111110110011110100001000000, 37'b1111111111111111101010101100100001110, 37'b0000000000000000000000000001001011001, 37'b0000000000000000111111110111011000110, 37'b1111111111111101100110000110101111011, 37'b0000000000000000110110011011100010011, 37'b0000000000000110100100110000000010000, 37'b0000000000000110110100101001111110000, 37'b0000000000000110001111111100011011111, 37'b0000000000000100111011011011100000011, 37'b0000000000000000000000001100011110111, 37'b0000000000000001110100111110000010000, 37'b0000000000001100100010010101111111110},
{37'b1111111111111111100110001011100101000, 37'b1111111111111100001100011110011011011, 37'b0000000000000110001110101101011101101, 37'b1111111111111110010110101010011001101, 37'b0000000000000001000111011101011000010, 37'b0000000000000010101011111001011111010, 37'b1111111111111111111111111111101010100, 37'b1111111111111011011010001010010000010, 37'b1111111111111110101000110001010010100, 37'b1111111111110110011000110111100010010, 37'b0000000000000111001010000010101100010, 37'b0000000000000000000011111000111001010, 37'b0000000000000110101101001000011101111, 37'b0000000000001010101110001101100110100, 37'b1111111111111110001000110011011110001, 37'b1111111111110010000100011101110100000, 37'b1111111111111110010101101010101100010, 37'b0000000000000111100001001011100111010, 37'b1111111111111011011110010111011111100, 37'b1111111111111100101010010111000001011, 37'b0000000000000000111100110110100101110, 37'b0000000000000000000001000000100110011, 37'b1111111111110111010001111011000101010, 37'b1111111111111100111100001001111110001, 37'b1111111111111111010111110010110100110, 37'b1111111111111110000011010000111101011, 37'b0000000000000001110010111110101111100, 37'b0000000000001011010000011111110100010, 37'b0000000000000011111011011010001101011, 37'b1111111111111111111111111010000100110, 37'b0000000000000001010010101011101101010, 37'b0000000000000000011100010011010010111},
{37'b0000000000000000101011011101010100000, 37'b0000000000000111010000100110110000000, 37'b0000000000000000000000000111100110100, 37'b0000000000000100101110100110110001000, 37'b0000000000001101010011001110100111000, 37'b1111111111111101010001001011101000011, 37'b1111111111111111111111111011111110011, 37'b1111111111111111010010101011000001111, 37'b0000000000000100101100000010101101010, 37'b1111111111111100111011111001010100110, 37'b1111111111111111111110101011101011110, 37'b0000000000000101010101010100100101111, 37'b0000000000000000001000101101100011010, 37'b0000000000000000011100000101111000000, 37'b1111111111100111100100010100100001100, 37'b1111111111111110101110101100010010110, 37'b0000000000000000000000000000011001010, 37'b0000000000000011001101100000000110000, 37'b1111111111111111111100100100001010000, 37'b0000000000000100110001110010100100101, 37'b1111111111111111111111110001010111110, 37'b1111111111111101001111000110100110111, 37'b1111111111110111000000100111111100110, 37'b0000000000000010000101111110101111001, 37'b0000000000000100100100110000010111110, 37'b1111111111101110010000001111110001100, 37'b1111111111111111111111110010100011100, 37'b0000000000000000000000001011101100101, 37'b0000000000001000101101001011010101100, 37'b1111111111110011001011011011101001000, 37'b0000000000000000000001110110010100010, 37'b1111111111111111111001110001100001100},
{37'b0000000000000000001001101010000010001, 37'b1111111111111010100100001111011111101, 37'b0000000000000000110111010001000101101, 37'b1111111111111111110000101101100111100, 37'b0000000000000000110101010100011010001, 37'b0000000000001000011101110001010100010, 37'b1111111111110100011001110111001101000, 37'b0000000000000000100011001110110010001, 37'b0000000000000110110001100101010101100, 37'b1111111111111010100110101100111100011, 37'b1111111111111111101000001110110011110, 37'b0000000000000000110010000100011111101, 37'b1111111111111111110110110110110001111, 37'b0000000000000010110111001010111011010, 37'b0000000000000001101101111100100110100, 37'b1111111111111111101110111110011111000, 37'b0000000000000001000100101011010110110, 37'b0000000000000000000000010011010100011, 37'b0000000000000000010110000111111011110, 37'b0000000000000110000100111111100110010, 37'b1111111111111111100011010001000111001, 37'b1111111111111000010000000000010011110, 37'b1111111111110110010100100111010101110, 37'b1111111111111100111001101010001110000, 37'b1111111111110110100011001001010111000, 37'b0000000000000011010101000001001000100, 37'b0000000000001001111110001101001010100, 37'b0000000000000101111001100001100111001, 37'b1111111111111111110101010101000101011, 37'b1111111111111010000010011100011001101, 37'b1111111111111011000001110011010011000, 37'b0000000000000000111101001011100100001},
{37'b0000000000000000110101001011001111010, 37'b1111111111111000010110111011001100101, 37'b1111111111111111101110101100110111001, 37'b0000000000000010011010000110010011000, 37'b1111111111111000010110000011000011001, 37'b0000000000000010101101110011101110111, 37'b1111111111111111111111111000001011010, 37'b1111111111111111111111110101011111101, 37'b1111111111111111111111111101101010001, 37'b0000000000000000000000001110010111101, 37'b0000000000000100001110101110101000000, 37'b1111111111111111101110010101111010010, 37'b0000000000000000001001111111000001110, 37'b0000000000000000000000010000100100010, 37'b0000000000000010000010011011000111000, 37'b1111111111111111101110101111101000100, 37'b0000000000000000000010110100101110000, 37'b1111111111111111111111010011111000110, 37'b1111111111111010110110001111100100111, 37'b1111111111110111111010001110000111100, 37'b1111111111111111111111011010001001000, 37'b1111111111110111011101010100011110100, 37'b1111111111111011001011100110111101001, 37'b1111111111111010000011010101101001011, 37'b0000000000001110001111111101010000100, 37'b0000000000000000010010000000100001000, 37'b1111111111111111010000110111100100011, 37'b0000000000000101000100111101011001011, 37'b0000000000001110010111000000000010010, 37'b0000000000000110010100010110101001110, 37'b1111111111101111000010000110000011000, 37'b1111111111111101000010000011010000001},
{37'b0000000000000110000000111001100001100, 37'b1111111111111111111111100110111100001, 37'b0000000000000100000001000011011101110, 37'b1111111111111111101011101010101011000, 37'b0000000000000111101111010111100100101, 37'b1111111111111101101101111110111110001, 37'b0000000000000001001000100001011111111, 37'b0000000000000110101100010001001101110, 37'b0000000000000100010010001101111110111, 37'b1111111111110111101001010001011110100, 37'b1111111111111111000000111111111000001, 37'b0000000000000001111101110100001011101, 37'b0000000000000001000110100111000101101, 37'b1111111111111111110001000010110100101, 37'b0000000000000001010110111100011100001, 37'b0000000000000000000000010001001111011, 37'b0000000000000101110011000100100110000, 37'b0000000000000000100011111010001110001, 37'b0000000000000101111111001011101110111, 37'b1111111111111110111100111011011011011, 37'b1111111111111101111101100111101001111, 37'b1111111111111110110011011001101101111, 37'b1111111111111111111111110000110111000, 37'b0000000000000100110101000110111110001, 37'b1111111111111100110000110010111101011, 37'b1111111111111111111001101001010000111, 37'b0000000000000000000000000000101010011, 37'b0000000000000000000000010000111111010, 37'b0000000000000000000000001000010000000, 37'b0000000000000100101011000111000011000, 37'b1111111111111010110111101000101111010, 37'b1111111111111111101000001110011111111},
{37'b1111111111111111111111010101110111010, 37'b1111111111111111100000011000111110010, 37'b1111111111111000100011110001100100110, 37'b0000000000000100100011010101101100001, 37'b0000000000000011100100100001000011010, 37'b1111111111111110001111110011010000111, 37'b1111111111111111111111110111101001011, 37'b1111111111111100010111101000101111001, 37'b0000000000000000000110111001001010111, 37'b1111111111111111111111101010101111000, 37'b1111111111111011001011011001011110110, 37'b1111111111111100000011110000110011001, 37'b0000000000000111101010100001111111001, 37'b0000000000000000000000000000101100010, 37'b1111111111111101111101001100000001011, 37'b1111111111111111111111111100100111110, 37'b0000000000000011011011001110000010110, 37'b1111111111111111111111110101100110100, 37'b1111111111111111111111111110110000110, 37'b1111111111111100100010110110100101011, 37'b0000000000000101000011111010011011011, 37'b0000000000000000000000000100011100001, 37'b0000000000000010011111111011111011110, 37'b1111111111111111100010101011110110101, 37'b0000000000000010100000110001000010000, 37'b0000000000000000000010010000100110010, 37'b0000000000000000000000000110110011011, 37'b0000000000000011110110100010000111000, 37'b1111111111111100111011010010110111111, 37'b1111111111111111010000110100111010010, 37'b0000000000000010100100011011001111000, 37'b1111111111111110010011100110010100010},
{37'b1111111111111111101110110111110011111, 37'b1111111111111011000100000001111100101, 37'b0000000000001001100000101010110011100, 37'b1111111111111110111101011111010010101, 37'b0000000000000011001001000111010101010, 37'b1111111111111011011011000011111001011, 37'b0000000000000000000000000100010100100, 37'b0000000000000000100011000000000010110, 37'b1111111111111000010101011110010000010, 37'b1111111111111111110010111010000110100, 37'b1111111111111110000001010001010011001, 37'b0000000000000000111011100100100101100, 37'b1111111111111010110000001111101100101, 37'b0000000000000010001101001101000001001, 37'b0000000000000011001111001000100101000, 37'b0000000000000001110000001101101110010, 37'b0000000000000001010111110110111001110, 37'b1111111111111111011001000011000110010, 37'b1111111111110100101010110101011000010, 37'b1111111111111111110010001101001110110, 37'b1111111111111111000101101110010111101, 37'b0000000000000010001111001100111010100, 37'b1111111111111110001110010000110110011, 37'b1111111111111111111111111111100001101, 37'b0000000000000011001010011101010000010, 37'b1111111111111111010001010110111111011, 37'b1111111111111111110001001101001001101, 37'b0000000000000110001110010110100101110, 37'b1111111111111001101000011100000010001, 37'b1111111111111011010001110000100110011, 37'b0000000000000101100111001111010000011, 37'b0000000000000000100100110001010011000},
{37'b0000000000000110111001010010011100101, 37'b0000000000000011001110001000101011011, 37'b0000000000000000000000110010001000010, 37'b1111111111111101011101001101110011111, 37'b1111111111111110101111101000110111010, 37'b1111111111111111111111001000110010001, 37'b0000000000000000000000000100100101010, 37'b1111111111111110111001001101101011000, 37'b1111111111111110000000110101000010110, 37'b1111111111111110000110101010101100101, 37'b0000000000000000000000010101010000111, 37'b0000000000000010100010001011100100110, 37'b0000000000000000000110100011000001000, 37'b0000000000000000110110001000001110010, 37'b1111111111111111010010010010000111100, 37'b0000000000000000000101111010000110001, 37'b1111111111111101100010111100110010101, 37'b0000000000000000000000100111000111110, 37'b1111111111111111101101111111110000001, 37'b1111111111111111111111011001101001110, 37'b0000000000000000000010011001011000011, 37'b0000000000000000111100110110110101000, 37'b0000000000000001100011100001100110111, 37'b0000000000000000000000000110000110001, 37'b0000000000000000000000010010001100000, 37'b1111111111110110001110110111100001100, 37'b1111111111111100110011111101001111011, 37'b0000000000000000000110110001000000101, 37'b0000000000000000010100111101001110001, 37'b0000000000000000000001010111000101111, 37'b1111111111111101001010101001011000000, 37'b0000000000000000010101111111111111100},
{37'b0000000000000011000000001000110100111, 37'b1111111111101111010010011001011100000, 37'b1111111111111111111111111001110100111, 37'b1111111111111110110010111110010000001, 37'b1111111111111100010001100010100110110, 37'b1111111111111111110110001011101111110, 37'b0000000000000000000000000010111101110, 37'b0000000000001000110000111100110111100, 37'b1111111111111111010011001000001101111, 37'b1111111111111111101001100000010101001, 37'b0000000000000001010100011111111100011, 37'b1111111111110101011011011101000001100, 37'b0000000000000000011000100100101001100, 37'b1111111111111000111111000001000001111, 37'b0000000000001011100011110001110001010, 37'b1111111111111111001010011110101000111, 37'b1111111111111100011000000110000000001, 37'b1111111111110111001111110111000010000, 37'b1111111111111111110101001110101111110, 37'b1111111111110100101011001101011100010, 37'b1111111111110011000010111000000001110, 37'b1111111111111111111111101101111111000, 37'b0000000000000000000000011101011101111, 37'b0000000000000000000000000100101101110, 37'b0000000000000011111001111000110011110, 37'b1111111111111111110001101111011101110, 37'b1111111111111011001110101001010100110, 37'b1111111111111110110101100100110000000, 37'b1111111111111111101000001000100011100, 37'b0000000000000000000000001110110111110, 37'b1111111111111111011111100010111010100, 37'b1111111111110100110011010000011111000}
};
localparam logic signed [36:0] bias [32] = '{
37'b0000000000000100001110011000101001100,
37'b0000000000000110101110110100001011011,
37'b0000000000000011001011101100000111010,
37'b0000000000000011010010001110011111000,
37'b1111111111100010101111001111010100100,
37'b1111111111111000110100010100111101111,
37'b0000000000001101101001000011110010010,
37'b1111111111110101110010011011001101000,
37'b1111111111111011010101000110101101100,
37'b0000000000010101100110001110110110100,
37'b0000000000000001101111001000111001011,
37'b0000000000000111000011010011101001010,
37'b1111111111101010111011001111001110100,
37'b1111111111110000111110110100101110010,
37'b0000000000001101010011001111000100110,
37'b0000000000010101111101111011111101100,
37'b1111111111111100001011000100011011101,
37'b0000000000001101100101101000011010000,
37'b0000000000000110110101101100111001110,
37'b0000000000001000000010010101110100000,
37'b0000000000001011010110111010110111000,
37'b0000000000000110101010001110001011001,
37'b0000000000000100010110001110101110000,
37'b0000000000000111011010111111110111110,
37'b1111111111111101010000100101010001110,
37'b1111111111111011100001111100001000001,
37'b1111111111111011000010000111100101000,
37'b1111111111110101110000100000101001000,
37'b0000000000000000011110011010011111110,
37'b1111111111111001011011011110100001100,
37'b0000000000000111000001101111010000100,
37'b1111111111111000011001110000001101011
};
endpackage