package softmax_exp_16_10;

localparam logic signed [15:0] exp_table [1023:0]= {
16'h00400,
16'h00AE0,
16'h01D8E,
16'h05058,
16'h0DA65,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h1FFFF,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00000,
16'h00001,
16'h00003,
16'h00007,
16'h00013,
16'h00033,
16'h0008B,
16'h00179
};
endpackage