// Width: 6
// NFRAC: 3
package dense_4_6_3;

localparam logic signed [5:0] weights [32][5] = '{ 
{6'b111111, 6'b000010, 6'b111101, 6'b000000, 6'b111111}, 
{6'b111011, 6'b111111, 6'b000011, 6'b111111, 6'b000000}, 
{6'b000010, 6'b000001, 6'b111111, 6'b111100, 6'b111110}, 
{6'b111100, 6'b111101, 6'b111111, 6'b000010, 6'b000001}, 
{6'b000000, 6'b000001, 6'b000001, 6'b111111, 6'b110111}, 
{6'b000010, 6'b111100, 6'b000001, 6'b111110, 6'b111110}, 
{6'b111100, 6'b000000, 6'b111111, 6'b000001, 6'b000000}, 
{6'b111111, 6'b000010, 6'b111100, 6'b000001, 6'b000001}, 
{6'b000001, 6'b111110, 6'b000000, 6'b111100, 6'b111110}, 
{6'b111111, 6'b111101, 6'b000001, 6'b000011, 6'b000000}, 
{6'b111110, 6'b111110, 6'b000000, 6'b000100, 6'b111101}, 
{6'b000001, 6'b000001, 6'b111101, 6'b111111, 6'b000000}, 
{6'b000000, 6'b000001, 6'b000000, 6'b111110, 6'b111011}, 
{6'b000001, 6'b000000, 6'b000011, 6'b111111, 6'b111100}, 
{6'b000000, 6'b111111, 6'b111101, 6'b111111, 6'b000100}, 
{6'b111100, 6'b111110, 6'b111110, 6'b000011, 6'b000000}, 
{6'b000010, 6'b111110, 6'b111110, 6'b111110, 6'b111111}, 
{6'b000001, 6'b111111, 6'b111100, 6'b111111, 6'b000000}, 
{6'b000010, 6'b000000, 6'b111110, 6'b000000, 6'b111100}, 
{6'b000001, 6'b111111, 6'b111110, 6'b000001, 6'b000000}, 
{6'b000000, 6'b111111, 6'b000010, 6'b111100, 6'b111111}, 
{6'b000000, 6'b000000, 6'b000011, 6'b111011, 6'b111011}, 
{6'b111111, 6'b000000, 6'b000001, 6'b111101, 6'b000100}, 
{6'b111111, 6'b000001, 6'b000010, 6'b000000, 6'b111011}, 
{6'b111110, 6'b000010, 6'b111110, 6'b000000, 6'b000011}, 
{6'b000000, 6'b000010, 6'b000000, 6'b111010, 6'b000100}, 
{6'b111100, 6'b111110, 6'b000001, 6'b000001, 6'b000001}, 
{6'b000000, 6'b000001, 6'b111111, 6'b111110, 6'b000000}, 
{6'b111111, 6'b000001, 6'b111011, 6'b000001, 6'b111110}, 
{6'b111111, 6'b000001, 6'b111110, 6'b111100, 6'b000100}, 
{6'b000011, 6'b000000, 6'b000010, 6'b111011, 6'b111101}, 
{6'b111111, 6'b111100, 6'b000010, 6'b000000, 6'b000001}
};

localparam logic signed [5:0] bias [5] = '{
6'b111111,  // -0.06223141402006149
6'b111111,  // -0.06270556896924973
6'b111111,  // -0.07014333456754684
6'b000000,  // 0.0820775106549263
6'b000001   // 0.2155742198228836
};
endpackage