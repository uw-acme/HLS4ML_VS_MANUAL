// Width: 21
// NFRAC: 10
package dense_2_21_10;

localparam logic signed [20:0] weights [64][32] = '{ 
{21'b000000000000100010011, 21'b000000000000000001000, 21'b111111111111100111101, 21'b111111111111111101010, 21'b000000000000100001011, 21'b000000000000000000000, 21'b111111111111101101100, 21'b111111111111111111111, 21'b111111111111011100111, 21'b000000000000001010001, 21'b000000000000000000000, 21'b111111111111111111010, 21'b111111111111111111111, 21'b111111111111100110011, 21'b111111111111111001100, 21'b111111111111011110011, 21'b000000000000000000000, 21'b111111111111111110010, 21'b111111111111100111100, 21'b111111111111101011101, 21'b000000000000000000000, 21'b000000000000000000000, 21'b111111111111111110111, 21'b111111111111111111101, 21'b000000000000000000000, 21'b000000000000001100110, 21'b000000000000110001011, 21'b000000000000010110011, 21'b111111111111111111111, 21'b000000000000000110011, 21'b111111111111001011100, 21'b000000000000000000000}, 
{21'b111111111111110011001, 21'b111111111111101100001, 21'b111111111111101110010, 21'b111111111111111000111, 21'b111111111111111111010, 21'b000000000000000101100, 21'b111111111111100011011, 21'b000000000000000000101, 21'b000000000000000000100, 21'b111111111111110111111, 21'b000000000000010011111, 21'b111111111111111010011, 21'b111111111111111000011, 21'b111111111111100100001, 21'b000000000000000000111, 21'b111111111111111001110, 21'b000000000000000001100, 21'b111111111111100111000, 21'b000000000000010101111, 21'b000000000000011101011, 21'b111111111111111011111, 21'b111111111111111111010, 21'b111111111111111111111, 21'b000000000000000011000, 21'b111111111111110110111, 21'b000000000000100011001, 21'b000000000000011111101, 21'b000000000000000001000, 21'b000000000000000011101, 21'b111111111111000001101, 21'b000000000000000000111, 21'b000000000000000000000}, 
{21'b000000000000001001010, 21'b111111111111110001010, 21'b111111111111101111011, 21'b111111111111111010101, 21'b111111111111110110000, 21'b111111111111110101000, 21'b111111111111101000010, 21'b000000000000000000100, 21'b111111111111101110101, 21'b000000000000000001001, 21'b000000000000000000010, 21'b111111111111110101101, 21'b000000000000001011100, 21'b111111111111110111101, 21'b111111111111111111110, 21'b111111111111111011010, 21'b000000000000000000101, 21'b000000000000001100001, 21'b000000000000000111100, 21'b000000000000011101011, 21'b000000000000000101010, 21'b111111111111110101001, 21'b000000000000000000000, 21'b000000000000000100011, 21'b111111111111111101101, 21'b000000000000011010110, 21'b000000000000010011000, 21'b000000000000001100011, 21'b111111111111111111111, 21'b111111111111101100100, 21'b111111111111111110010, 21'b000000000000001100101}, 
{21'b000000000000010001101, 21'b000000000000000010011, 21'b000000000000000110110, 21'b111111111111111110110, 21'b111111111110111110110, 21'b000000000000000000000, 21'b000000000000000000000, 21'b000000000000011100111, 21'b000000000000011111000, 21'b111111111111111110010, 21'b111111111111111111111, 21'b000000000000000000000, 21'b000000000000000000000, 21'b000000000000000000101, 21'b111111111111111101101, 21'b000000000000011011011, 21'b000000000000000000000, 21'b111111111111111100110, 21'b111111111111111111111, 21'b111111111111101001011, 21'b111111111111111000001, 21'b000000000000000110010, 21'b111111111111110111111, 21'b111111111111111111111, 21'b000000000000000000011, 21'b111111111111111001100, 21'b000000000000001001010, 21'b111111111111111111111, 21'b111111111111111111111, 21'b111111111111111111111, 21'b111111111111100100011, 21'b000000000000100111101}, 
{21'b111111111110101000101, 21'b111111111111111100110, 21'b111111111111111111011, 21'b000000000000000000101, 21'b111111111111111100101, 21'b000000000000000000110, 21'b111111111111111001101, 21'b111111111111101100110, 21'b000000000000000110111, 21'b111111111111111101011, 21'b111111111111111110010, 21'b111111111111111111111, 21'b111111111111111111111, 21'b000000000000011010111, 21'b000000000000000000000, 21'b000000000000101010000, 21'b111111111111111111111, 21'b000000000000011011111, 21'b111111111111001100110, 21'b000000000000000000000, 21'b111111111111110001101, 21'b000000000000010101100, 21'b000000000000100001000, 21'b000000000000000000000, 21'b000000000000000101110, 21'b000000000000010100110, 21'b000000000000011110100, 21'b000000000000000010001, 21'b111111111111111111011, 21'b111111111111111111111, 21'b111111111111111110001, 21'b000000000000011100111}, 
{21'b000000000000000111011, 21'b111111111111111111111, 21'b000000000000010011000, 21'b111111111110101100111, 21'b111111111101001111101, 21'b111111111111010011001, 21'b000000000000101101010, 21'b111111111110110000010, 21'b111111111111111111111, 21'b111111111110101001010, 21'b111111111110111111110, 21'b111111111111010100010, 21'b000000000000101101001, 21'b111111111111111111111, 21'b111111111111111110000, 21'b000000000000000000000, 21'b111111111111111111111, 21'b111111111111111111111, 21'b111111111111101111000, 21'b111111111111111111111, 21'b111111111111000001011, 21'b000000000000000000000, 21'b000000000000010111110, 21'b111111111111111111111, 21'b000000000000000010110, 21'b000000000000100010010, 21'b000000000000000110100, 21'b111111111111111111111, 21'b111111111111111111111, 21'b000000000000011010010, 21'b111111111111111011101, 21'b000000000000011001101}, 
{21'b111111111111111011011, 21'b111111111111101011110, 21'b111111111111100001000, 21'b111111111111111001111, 21'b111111111111011011000, 21'b000000000000001000011, 21'b111111111111101000111, 21'b111111111111101101110, 21'b111111111111001010111, 21'b000000000000000110001, 21'b111111111111111111010, 21'b111111111111101011101, 21'b000000000000001111001, 21'b111111111111111110101, 21'b111111111111111010101, 21'b111111111110111001001, 21'b111111111111111111111, 21'b000000000000001010110, 21'b000000000000011000100, 21'b111111111111101011001, 21'b111111111111101100110, 21'b111111111111110111111, 21'b111111111111111111110, 21'b000000000000000011100, 21'b111111111111111010001, 21'b111111111110101101000, 21'b111111111111011110000, 21'b111111111111111010001, 21'b000000000000000000101, 21'b111111111111111101010, 21'b000000000000000011111, 21'b111111111111111111111}, 
{21'b111111111111101100010, 21'b111111111111110100011, 21'b111111111111110101110, 21'b111111111111100001101, 21'b111111111111110001001, 21'b111111111111111111111, 21'b000000000000001101010, 21'b111111111111110101111, 21'b000000000000011001101, 21'b000000000000000000000, 21'b000000000000000000000, 21'b111111111111111111111, 21'b000000000000011100000, 21'b000000000000000000000, 21'b111111111111111111111, 21'b111111111111110110111, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111111111111, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111111111111, 21'b000000000000000101101, 21'b111111111111101000111, 21'b000000000000000001110, 21'b111111111111111111111, 21'b111111111111110110110, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111111111111}, 
{21'b111111111111000010111, 21'b111111111111111000101, 21'b111111111111001111010, 21'b000000000000001111101, 21'b000000000000111110010, 21'b111111111111111111111, 21'b111111111111111100010, 21'b000000000000011110100, 21'b111111111111000111110, 21'b111111111111111010000, 21'b000000000000000000000, 21'b111111111111100110001, 21'b111111111111111111111, 21'b000000000000001001101, 21'b111111111111100111100, 21'b000000000001100000100, 21'b111111111111111110111, 21'b000000000000000101111, 21'b000000000000011010100, 21'b000000000000011111010, 21'b000000000000000000000, 21'b111111111111010101000, 21'b000000000000000000000, 21'b000000000000110100101, 21'b111111111111101000110, 21'b000000000001011001010, 21'b111111111111101100111, 21'b111111111111100101111, 21'b111111111111000011100, 21'b111111111111000100100, 21'b000000000000000000000, 21'b000000000000000110110}, 
{21'b000000000000000000000, 21'b111111111111111110000, 21'b111111111111110110100, 21'b000000000000000000000, 21'b000000000000100111011, 21'b111111111111111101011, 21'b111111111111110111110, 21'b000000000000001011110, 21'b000000000000001100111, 21'b000000000000000000011, 21'b111111111111111110111, 21'b111111111111111111111, 21'b111111111111111111111, 21'b111111111111110001011, 21'b111111111111111111111, 21'b000000000000000000000, 21'b000000000000000000000, 21'b111111111111111111010, 21'b000000000000000000010, 21'b000000000000001010110, 21'b000000000000000010011, 21'b111111111111111111111, 21'b000000000000000000000, 21'b000000000000000000111, 21'b000000000000000100111, 21'b111111111111101111000, 21'b000000000000001000101, 21'b000000000000011111110, 21'b111111111111111111111, 21'b000000000000000000110, 21'b000000000000000110010, 21'b000000000000001000111}, 
{21'b000000000000001100010, 21'b000000000000000000000, 21'b111111111111110010110, 21'b111111111111011111111, 21'b111111111110011010010, 21'b000000000000010001000, 21'b000000000000000000000, 21'b111111111110010110000, 21'b000000000000000100101, 21'b111111111111111111111, 21'b000000000000000000011, 21'b111111111111111111110, 21'b000000000000000001010, 21'b000000000000000000000, 21'b111111111111111101100, 21'b111111111111001111001, 21'b111111111111111111111, 21'b000000000000011100001, 21'b000000000000010000001, 21'b000000000000011000011, 21'b111111111111000111101, 21'b111111111111010010011, 21'b000000000000001111010, 21'b111111111111111011100, 21'b111111111111111010000, 21'b000000000000101101111, 21'b111111111111110011101, 21'b111111111111111111111, 21'b111111111111111111111, 21'b000000000000011011000, 21'b111111111111111111111, 21'b000000000000000000110}, 
{21'b111111111111100110101, 21'b111111111111000000111, 21'b000000000000000000000, 21'b111111111111111111101, 21'b000000000000101010100, 21'b111111111111011101100, 21'b111111111111100011101, 21'b000000000000001110110, 21'b111111111111111111111, 21'b000000000000010011000, 21'b000000000000001001011, 21'b111111111111110110010, 21'b000000000000000000000, 21'b000000000000000001110, 21'b111111111111111101010, 21'b111111111111011111100, 21'b000000000000010110011, 21'b000000000000000011101, 21'b000000000000100110000, 21'b000000000000001011000, 21'b000000000000000000000, 21'b111111111111111011001, 21'b000000000000010000001, 21'b111111111111110100111, 21'b111111111111011000100, 21'b111111111111111111001, 21'b000000000000010111101, 21'b111111111111111111111, 21'b000000000000000001000, 21'b111111111111110011111, 21'b000000000000010001100, 21'b000000000000100011010}, 
{21'b000000000000000001111, 21'b000000000000000000000, 21'b000000000000011100000, 21'b000000000000000001000, 21'b111111111111111010110, 21'b000000000000010111000, 21'b000000000000001011110, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111101110000, 21'b111111111111111001000, 21'b111111111111101010100, 21'b111111111111111111111, 21'b000000000000000110011, 21'b111111111111110111001, 21'b000000000001101011111, 21'b000000000000000000000, 21'b111111111111110011111, 21'b111111111111100111110, 21'b111111111111111110010, 21'b000000000000011001011, 21'b000000000000010000011, 21'b000000000000000000000, 21'b111111111111111111101, 21'b000000000000011100000, 21'b000000000000100010010, 21'b000000000000111111011, 21'b000000000000000001010, 21'b000000000000000000000, 21'b000000000000000000000, 21'b111111111111111110011, 21'b111111111111110110110}, 
{21'b111111111111101100000, 21'b000000000000000110001, 21'b000000000000000101000, 21'b111111111111100000010, 21'b111111111111011101100, 21'b000000000000111100000, 21'b000000000000000110010, 21'b000000000000000000000, 21'b111111111111101011011, 21'b111111111111110100101, 21'b000000000000010000100, 21'b000000000000001001000, 21'b000000000000000000000, 21'b111111111111110101111, 21'b000000000000100100100, 21'b111111111111111111111, 21'b111111111111111110010, 21'b000000000000000000000, 21'b000000000000000001101, 21'b111111111111111010000, 21'b000000000000001010000, 21'b000000000000000010000, 21'b000000000000001110100, 21'b111111111111111111111, 21'b000000000000000000011, 21'b000000000001010100001, 21'b111111111111111000110, 21'b111111111111111101000, 21'b111111111111111111111, 21'b111111111111110010000, 21'b111111111111111010110, 21'b000000000000010110100}, 
{21'b000000000000000111100, 21'b000000000000001001011, 21'b000000000000101001110, 21'b111111111111111010111, 21'b000000000000001100111, 21'b000000000000101100111, 21'b000000000000000000000, 21'b111111111111111100001, 21'b000000000000001111000, 21'b111111111111110001011, 21'b111111111111111111111, 21'b111111111111110000101, 21'b000000000000000000000, 21'b000000000000110010010, 21'b111111111111111101101, 21'b000000000000000000001, 21'b000000000000011110001, 21'b000000000000000000000, 21'b000000000000000000011, 21'b111111111111010111111, 21'b111111111111100000100, 21'b111111111111111011011, 21'b111111111111111111111, 21'b111111111111101101010, 21'b111111111111111011011, 21'b111111111111110101011, 21'b111111111111100110110, 21'b111111111111100100110, 21'b000000000000000011110, 21'b000000000000001110010, 21'b111111111111001101001, 21'b000000000000000000011}, 
{21'b111111111111011001110, 21'b000000000000000000000, 21'b111111111111111110000, 21'b111111111111111001101, 21'b111111111111111111111, 21'b000000000000010001000, 21'b111111111111110110000, 21'b000000000000100010101, 21'b111111111111010001100, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111111111111, 21'b000000000000000000000, 21'b000000000000000000000, 21'b111111111111111111100, 21'b111111111111110100011, 21'b000000000000001010001, 21'b000000000000010111011, 21'b111111111111111110110, 21'b111111111111011111110, 21'b111111111111111000011, 21'b000000000000001110010, 21'b000000000000001000000, 21'b000000000000000000000, 21'b000000000000000000011, 21'b000000000000001010011, 21'b111111111111100001010, 21'b000000000000000000000, 21'b111111111111111111111, 21'b000000000000000000011, 21'b000000000000000000000, 21'b111111111111101111111}, 
{21'b111111111111010100111, 21'b111111111111111111010, 21'b111111111111111111100, 21'b111111111111111101110, 21'b111111111111111111011, 21'b000000000000001101100, 21'b000000000000000000110, 21'b000000000000000100011, 21'b000000000000000100111, 21'b000000000000001000000, 21'b000000000000001010000, 21'b000000000000010100101, 21'b000000000000000011011, 21'b111111111111110011100, 21'b000000000000000000000, 21'b000000000000110000110, 21'b000000000000000000000, 21'b000000000000000000001, 21'b111111111111111111101, 21'b000000000000001110000, 21'b000000000000010010001, 21'b000000000000000011111, 21'b000000000000000101010, 21'b111111111111111100001, 21'b111111111111111011111, 21'b000000000000000011011, 21'b111111111111110111011, 21'b111111111111101111110, 21'b000000000000011010110, 21'b111111111111111100000, 21'b000000000000000100000, 21'b111111111111100111111}, 
{21'b000000000000000000000, 21'b111111111111111111111, 21'b000000000000000100110, 21'b000000000000000000000, 21'b000000000001110100000, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111111111111, 21'b000000000000001110000, 21'b111111111111110110011, 21'b000000000000000000000, 21'b000000000000000000000, 21'b000000000000000000001, 21'b000000000000010000100, 21'b000000000000000000000, 21'b111111111111101101011, 21'b111111111111111111111, 21'b111111111111110111011, 21'b000000000000101001111, 21'b000000000000000000000, 21'b111111111111111111111, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111111111111, 21'b000000000000000000000, 21'b000000000000001000101, 21'b000000000000000000000, 21'b000000000000000000000, 21'b111111111111111111111, 21'b111111111111111111111, 21'b000000000000000000000, 21'b000000000000000101010}, 
{21'b111111111111111111100, 21'b000000000000000011101, 21'b111111111111111111111, 21'b000000000000000110001, 21'b111111111111111010010, 21'b111111111111110000101, 21'b111111111111111000000, 21'b000000000000100011100, 21'b000000000000000000000, 21'b000000000000001100011, 21'b111111111111111110100, 21'b000000000000001000010, 21'b111111111111111011110, 21'b111111111111101011110, 21'b111111111111100111100, 21'b000000000000000001101, 21'b111111111111111111111, 21'b111111111111111011100, 21'b000000000000000000000, 21'b000000000000000000000, 21'b111111111111111111111, 21'b000000000000001001101, 21'b000000000000000100100, 21'b111111111111101111111, 21'b000000000000001110010, 21'b111111111111101010111, 21'b000000000000000000010, 21'b000000000000000000000, 21'b111111111111101010100, 21'b000000000000000000000, 21'b000000000000000101110, 21'b111111111111111100000}, 
{21'b111111111111111110100, 21'b111111111111110011010, 21'b000000000000000000000, 21'b111111111111111000010, 21'b000000000000011011101, 21'b111111111111111111111, 21'b111111111111111101010, 21'b000000000000001101101, 21'b111111111111001101111, 21'b000000000000000000000, 21'b111111111111111011000, 21'b111111111111111111101, 21'b000000000000101100111, 21'b000000000000011101010, 21'b111111111111110011010, 21'b111111111111111101010, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111111111111, 21'b000000000000000000000, 21'b000000000000000000000, 21'b111111111111101110100, 21'b111111111111110000110, 21'b000000000000010000110, 21'b000000000000000000000, 21'b111111111111101110011, 21'b000000000000000011001, 21'b111111111111110101101, 21'b111111111111111011101, 21'b000000000000010001011, 21'b000000000000000000000, 21'b111111111111100000010}, 
{21'b000000000001010001001, 21'b000000000000101011110, 21'b111111111111100000000, 21'b000000000000000000011, 21'b111111111111010011101, 21'b000000000000000000000, 21'b000000000000011100100, 21'b000000000000000011111, 21'b000000000000011100101, 21'b111111111111111111111, 21'b111111111111101100001, 21'b111111111111110101111, 21'b000000000000010010001, 21'b000000000000000011100, 21'b111111111111110011011, 21'b000000000000010000110, 21'b000000000001000100100, 21'b111111111111101111010, 21'b111111111111011010000, 21'b000000000000000000000, 21'b111111111111111100010, 21'b111111111111101001011, 21'b111111111111111110011, 21'b111111111111111111110, 21'b000000000000001011000, 21'b111111111111010001110, 21'b000000000000001011011, 21'b111111111111111111110, 21'b000000000000000000000, 21'b000000000000001101111, 21'b111111111111111100010, 21'b000000000000000111101}, 
{21'b111111111111110100001, 21'b111111111111100111011, 21'b111111111111111011010, 21'b111111111111101010100, 21'b111111111111111101110, 21'b000000000000000110010, 21'b000000000000000000000, 21'b111111111111111110100, 21'b000000000000000100110, 21'b111111111111111111100, 21'b000000000000000000000, 21'b111111111111100100001, 21'b000000000000001101000, 21'b000000000000001010010, 21'b111111111111110010111, 21'b000000000000111000110, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111111111011, 21'b000000000000000000000, 21'b000000000000101000011, 21'b111111111111000011110, 21'b111111111111110010001, 21'b111111111111111000110, 21'b111111111111111101100, 21'b000000000000011001001, 21'b111111111111111001010, 21'b000000000000000010010, 21'b000000000000111101111, 21'b111111111110111110011, 21'b111111111111010001000, 21'b000000000000000010110}, 
{21'b000000000000000010001, 21'b111111111111111000011, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111110100011111, 21'b111111111110110010011, 21'b000000000000000000001, 21'b111111111111111111111, 21'b111111111111011110000, 21'b000000000000000011001, 21'b000000000000000000000, 21'b111111111111111100011, 21'b000000000000000000000, 21'b111111111111111000100, 21'b111111111111111001010, 21'b111111111111110111001, 21'b111111111111101101001, 21'b000000000000100100001, 21'b000000000000000000000, 21'b000000000000000101111, 21'b111111111111111111111, 21'b111111111111110110111, 21'b000000000000000000000, 21'b111111111111110100111, 21'b000000000000011100000, 21'b111111111110110000010, 21'b000000000000011100001, 21'b111111111111111111111, 21'b111111111111111111011, 21'b000000000000011001100, 21'b111111111111111111111, 21'b000000000000011110001}, 
{21'b111111111111111111111, 21'b000000000000000000101, 21'b111111111111111010011, 21'b000000000000001001100, 21'b000000000000000111000, 21'b111111111111010100001, 21'b000000000000000000000, 21'b000000000000001000001, 21'b000000000001001010001, 21'b111111111111111110110, 21'b000000000000000000000, 21'b000000000000000111001, 21'b000000000000101101111, 21'b111111111111111011111, 21'b000000000000000001110, 21'b000000000000001100111, 21'b111111111111111111111, 21'b000000000000000011100, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111011100111, 21'b000000000000000100111, 21'b000000000000001000111, 21'b000000000000000010111, 21'b111111111111111111111, 21'b000000000000011011111, 21'b000000000000000000100, 21'b000000000000010000001, 21'b111111111111001010100, 21'b000000000000001101001, 21'b000000000000110010101, 21'b000000000000000000101}, 
{21'b111111111111010011000, 21'b000000000000011011000, 21'b111111111111011110101, 21'b000000000000001111101, 21'b111111111111110010100, 21'b000000000000000000000, 21'b000000000000111111101, 21'b111111111111100010001, 21'b111111111111011010101, 21'b000000000000010101111, 21'b111111111111100011011, 21'b111111111111111100111, 21'b111111111111111111111, 21'b000000000000101100000, 21'b111111111111111111110, 21'b111111111111011001011, 21'b111111111111111111111, 21'b000000000000111000011, 21'b111111111111000011101, 21'b111111111111111100111, 21'b000000000000101000100, 21'b111111111111010001100, 21'b000000000000000110110, 21'b111111111111111110000, 21'b000000000000100010101, 21'b111111111110111110111, 21'b111111111111010001100, 21'b111111111111100110111, 21'b111111111111111111111, 21'b000000000000001101010, 21'b000000000000000011001, 21'b000000000000010110110}, 
{21'b111111111111110100011, 21'b000000000000000110101, 21'b111111111111111111111, 21'b000000000000010011001, 21'b111111111111111011001, 21'b000000000000011101000, 21'b000000000000000000010, 21'b111111111111111110100, 21'b111111111111111111101, 21'b000000000000000000001, 21'b000000000000000000000, 21'b111111111111111111111, 21'b111111111111111111110, 21'b000000000001000010100, 21'b000000000000000001100, 21'b000000000000011000001, 21'b000000000000000000000, 21'b111111111111100100111, 21'b111111111111110110001, 21'b111111111111111111111, 21'b111111111111111101111, 21'b000000000000000101011, 21'b111111111111111111111, 21'b111111111111101000010, 21'b111111111111111111111, 21'b000000000000100101110, 21'b000000000000100111101, 21'b111111111111111111111, 21'b111111111111111101111, 21'b000000000000000000000, 21'b111111111111111111111, 21'b111111111111110011101}, 
{21'b111111111111110101101, 21'b000000000000000000000, 21'b000000000000100010111, 21'b000000000000000000000, 21'b000000000000000000000, 21'b111111111111110001011, 21'b000000000000000000000, 21'b111111111110010001011, 21'b000000000000011011100, 21'b000000000000000001110, 21'b000000000000000011011, 21'b111111111111010001111, 21'b000000000000000000011, 21'b111111111111101110011, 21'b111111111111111011110, 21'b000000000000000000000, 21'b000000000000000010100, 21'b000000000000000000000, 21'b000000000000001110011, 21'b000000000000000000000, 21'b111111111111111110110, 21'b000000000000101010001, 21'b000000000000110000001, 21'b111111111111100011101, 21'b111111111111101101110, 21'b000000000000011111111, 21'b111111111111011000111, 21'b000000000000000011110, 21'b111111111111111111111, 21'b111111111111111111111, 21'b111111111111111111111, 21'b000000000000010111100}, 
{21'b111111111111110001011, 21'b111111111111111111111, 21'b111111111111100001011, 21'b111111111111100110001, 21'b111111111111111110001, 21'b111111111111101110101, 21'b000000000000000000000, 21'b000000000000001011101, 21'b111111111111100001010, 21'b111111111111110101010, 21'b111111111111111001101, 21'b000000000000000000000, 21'b000000000000000011100, 21'b111111111111111110101, 21'b111111111111111000001, 21'b000000000000001100001, 21'b000000000000011100100, 21'b000000000000010000110, 21'b111111111111101111010, 21'b000000000000000110001, 21'b111111111111111110011, 21'b111111111111111100010, 21'b000000000000000010111, 21'b000000000000000010000, 21'b111111111111110111000, 21'b000000000000001011011, 21'b111111111111110100011, 21'b000000000000000111101, 21'b111111111111111111111, 21'b111111111111011010001, 21'b111111111111111100101, 21'b000000000000011100110}, 
{21'b111111111111111100100, 21'b111111111111110101011, 21'b000000000000001001110, 21'b000000000000100000011, 21'b000000000000001010110, 21'b000000000000001010100, 21'b000000000000000101111, 21'b111111111111100110001, 21'b111111111111100101101, 21'b000000000000001000110, 21'b000000000000000001100, 21'b000000000000000101100, 21'b000000000000000010110, 21'b000000000000000000101, 21'b000000000000011010010, 21'b000000000000000000111, 21'b111111111111111001000, 21'b000000000000001101001, 21'b111111111111111100001, 21'b111111111111111011011, 21'b000000000000001110000, 21'b111111111111110000001, 21'b111111111111111100100, 21'b000000000000010000010, 21'b000000000000000010110, 21'b111111111111110010010, 21'b111111111111100110101, 21'b111111111111111110011, 21'b111111111111011100010, 21'b000000000000000111101, 21'b000000000000001101000, 21'b000000000000000000001}, 
{21'b111111111111111110010, 21'b111111111111111101011, 21'b111111111111111110011, 21'b111111111111111011100, 21'b111111111111101111001, 21'b111111111111101110000, 21'b000000000000001000000, 21'b000000000000000001000, 21'b111111111111101000101, 21'b000000000000010101011, 21'b111111111111111101010, 21'b111111111111111111111, 21'b111111111111110001111, 21'b000000000000000000101, 21'b000000000000000011110, 21'b111111111111111001010, 21'b111111111111111101111, 21'b111111111111111010101, 21'b111111111111110101101, 21'b000000000000000000000, 21'b111111111111101110000, 21'b000000000000001101000, 21'b111111111111100100111, 21'b000000000000000000101, 21'b000000000000000101010, 21'b000000000000001111110, 21'b000000000000000011011, 21'b000000000000000000110, 21'b000000000000100101011, 21'b000000000000000110100, 21'b000000000000000000000, 21'b000000000000001010101}, 
{21'b111111111111111101100, 21'b000000000000100000010, 21'b111111111111111111111, 21'b111111111111111011110, 21'b111111111111100100101, 21'b111111111111110110011, 21'b000000000000110100101, 21'b111111111110100111110, 21'b111111111111010011010, 21'b111111111111100110011, 21'b111111111111100011111, 21'b111111111111011111100, 21'b111111111111111111111, 21'b000000000000111101111, 21'b111111111111111100101, 21'b000000000000000000000, 21'b111111111111100100111, 21'b000000000000111001000, 21'b111111111111001011001, 21'b000000000000000000000, 21'b111111111111111111111, 21'b111111111111010100111, 21'b000000000000000000000, 21'b111111111111111111111, 21'b000000000000000111001, 21'b111111111111111000101, 21'b111111111111101101000, 21'b111111111111111111111, 21'b000000000000010110010, 21'b000000000000000000011, 21'b111111111111110101101, 21'b000000000000000000000}, 
{21'b000000000000101111000, 21'b111111111111110001101, 21'b000000000000010000111, 21'b111111111111111011110, 21'b000000000000001001110, 21'b111111111111111111100, 21'b111111111111111111101, 21'b111111111111110100000, 21'b000000000000000000000, 21'b000000000000001011110, 21'b111111111111111111111, 21'b111111111111111000011, 21'b111111111111111111111, 21'b000000000000011101010, 21'b000000000000000010011, 21'b000000000000000101001, 21'b000000000000000011000, 21'b111111111111111100111, 21'b000000000000000010100, 21'b000000000000000000000, 21'b111111111111111110110, 21'b111111111111111111111, 21'b111111111111011000111, 21'b111111111111111111111, 21'b000000000000000111011, 21'b111111111111110001000, 21'b111111111111101110101, 21'b111111111111111111111, 21'b111111111111111111111, 21'b000000000001000111011, 21'b111111111111011011011, 21'b111111111111110001001}, 
{21'b111111111111111010010, 21'b111111111111110010110, 21'b111111111111110111101, 21'b000000000000000100101, 21'b000000000000010001110, 21'b111111111111101111011, 21'b111111111111111111110, 21'b111111111111100011110, 21'b000000000000000111110, 21'b000000000000010001011, 21'b111111111111100100101, 21'b111111111111011111101, 21'b000000000000000011000, 21'b111111111110101000100, 21'b111111111111110110010, 21'b111111111111110000001, 21'b111111111111100110101, 21'b111111111111111111111, 21'b000000000000010001001, 21'b000000000000000000000, 21'b111111111111111010001, 21'b111111111111111010010, 21'b000000000000000000000, 21'b000000000000000000000, 21'b111111111111111000011, 21'b111111111110011111011, 21'b111111111110111000111, 21'b111111111111011101000, 21'b000000000000000111001, 21'b000000000000011010011, 21'b111111111111111111111, 21'b000000000000011110110}, 
{21'b111111111111110100001, 21'b111111111111100100100, 21'b000000000000010100111, 21'b000000000000001001100, 21'b000000000000000101100, 21'b111111111111110100001, 21'b111111111111111011110, 21'b000000000000001100100, 21'b000000000001000100111, 21'b111111111111101010000, 21'b111111111111111111111, 21'b111111111111111111111, 21'b000000000000001111000, 21'b111111111111111000111, 21'b111111111111111101101, 21'b111111111111111101110, 21'b111111111111110011001, 21'b111111111111111111111, 21'b000000000000000000000, 21'b000000000000011101000, 21'b111111111111101110111, 21'b111111111111111111100, 21'b000000000000010000011, 21'b111111111111111110101, 21'b000000000000000000000, 21'b000000000001000011010, 21'b000000000000101001100, 21'b000000000000000000011, 21'b000000000000000000000, 21'b111111111111001010001, 21'b111111111111110111010, 21'b111111111111111111111}, 
{21'b000000000000000001111, 21'b000000000000000110001, 21'b111111111111111110001, 21'b000000000000000000000, 21'b000000000000011101100, 21'b111111111111000010001, 21'b000000000000000000000, 21'b111111111111110011110, 21'b000000000000010111110, 21'b000000000000000000000, 21'b111111111111111101101, 21'b000000000000000000000, 21'b000000000000000000000, 21'b111111111111111111111, 21'b000000000000000000101, 21'b111111111111110010001, 21'b000000000000100001001, 21'b111111111111111111010, 21'b111111111111111110000, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111111111000, 21'b000000000000000000000, 21'b111111111111111111111, 21'b000000000000000001101, 21'b111111111111010111011, 21'b000000000000000110100, 21'b000000000000010111011, 21'b111111111111111111100, 21'b000000000000001100000, 21'b111111111111111111111, 21'b000000000000001001100}, 
{21'b111111111111100110001, 21'b000000000000000001001, 21'b111111111111000010010, 21'b000000000000000000111, 21'b111111111111111001100, 21'b111111111111111010111, 21'b111111111111111111110, 21'b111111111111110100010, 21'b111111111111111011011, 21'b111111111111110111101, 21'b000000000000000110000, 21'b000000000000000011011, 21'b111111111111101001010, 21'b000000000000000000000, 21'b111111111111111111110, 21'b111111111111111110111, 21'b000000000000001001000, 21'b111111111111111101011, 21'b111111111111111100011, 21'b111111111111111100010, 21'b111111111111111111111, 21'b000000000000100010101, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111111110110, 21'b000000000000101000100, 21'b000000000000011000001, 21'b000000000000000100010, 21'b111111111111110011101, 21'b111111111111111110101, 21'b000000000000001000010, 21'b000000000000000111010}, 
{21'b000000000000000100010, 21'b000000000000000101000, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111000100000, 21'b000000000000000101100, 21'b000000000000000011001, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111101010010, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111101011011, 21'b000000000000000000000, 21'b000000000000000000000, 21'b000000000000000000000, 21'b000000000000000000000, 21'b111111111111010010011, 21'b000000000000000001001, 21'b111111111111111111111, 21'b111111111111111111111, 21'b000000000000000000000, 21'b000000000000010000100, 21'b111111111111111111111, 21'b000000000000000000000, 21'b000000000000111010010, 21'b000000000000101011100, 21'b000000000000000000000, 21'b000000000000000000000, 21'b111111111111100010000, 21'b000000000000000000000, 21'b111111111111111111111}, 
{21'b000000000000001001101, 21'b000000000000000110110, 21'b000000000000100000011, 21'b111111111111100000001, 21'b000000000000010000111, 21'b000000000000001111001, 21'b000000000000000000110, 21'b000000000000011000100, 21'b000000000000000001100, 21'b111111111111111110011, 21'b000000000000000100110, 21'b000000000000000000101, 21'b111111111111111111111, 21'b000000000000001111011, 21'b111111111111111111010, 21'b111111111111111010111, 21'b000000000000000000000, 21'b000000000000000100000, 21'b111111111111111001110, 21'b000000000000001100101, 21'b000000000000000100001, 21'b111111111110110101101, 21'b111111111111110001010, 21'b000000000000001011101, 21'b111111111111111111111, 21'b111111111110111111010, 21'b111111111111101111110, 21'b111111111111111101000, 21'b111111111111111111111, 21'b111111111111111000101, 21'b000000000000000000000, 21'b111111111111111010111}, 
{21'b000000000000000000001, 21'b111111111111111111111, 21'b111111111111110100010, 21'b111111111111101010011, 21'b000000000000000101010, 21'b000000000000000000000, 21'b000000000000001100001, 21'b111111111111111111010, 21'b000000000000011111111, 21'b111111111111111111011, 21'b000000000000000000000, 21'b111111111111010100000, 21'b111111111111111111111, 21'b000000000000010000000, 21'b111111111111111111111, 21'b111111111111011110101, 21'b000000000000000000000, 21'b111111111111111110100, 21'b000000000000100001101, 21'b111111111111111111111, 21'b111111111111001000000, 21'b111111111111111111111, 21'b000000000000100001000, 21'b111111111111111111111, 21'b111111111111111111111, 21'b000000000000010001110, 21'b111111111111110011111, 21'b000000000000001000110, 21'b000000000000000000000, 21'b111111111111100110001, 21'b000000000000000000000, 21'b000000000000000000010}, 
{21'b111111111111100100010, 21'b000000000000000000001, 21'b000000000000000000000, 21'b111111111111111111001, 21'b000000000000111111011, 21'b111111111111110000000, 21'b111111111111111111010, 21'b111111111111111111000, 21'b111111111111111010010, 21'b111111111111111001100, 21'b000000000000001000010, 21'b000000000000010001000, 21'b111111111111111011010, 21'b000000000000011111111, 21'b000000000000000000000, 21'b111111111111111111111, 21'b111111111111011011101, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111110101110, 21'b000000000000000000010, 21'b000000000000000100110, 21'b000000000000000001101, 21'b111111111111111110110, 21'b111111111111111001011, 21'b111111111111100110000, 21'b111111111111011010001, 21'b000000000000000000000, 21'b111111111111110001100, 21'b000000000000000101000, 21'b111111111111111111111, 21'b000000000000001001101}, 
{21'b111111111111001011000, 21'b111111111111101011111, 21'b111111111111101100000, 21'b000000000000000000000, 21'b000000000001001001000, 21'b111111111111100011100, 21'b000000000000000000000, 21'b111111111111111001000, 21'b111111111111001011100, 21'b000000000000010001101, 21'b111111111111111111111, 21'b000000000001001000100, 21'b000000000000000000000, 21'b111111111111111001111, 21'b111111111111111111111, 21'b000000000000000100000, 21'b111111111111111101100, 21'b000000000000000000000, 21'b111111111111111010000, 21'b000000000000111111011, 21'b000000000000000100111, 21'b111111111111111010101, 21'b000000000000001110000, 21'b111111111111111111111, 21'b111111111111111111111, 21'b111111111111110011100, 21'b111111111111111010000, 21'b111111111111000100000, 21'b111111111111101101100, 21'b111111111111111111111, 21'b111111111111111111110, 21'b111111111111111000011}, 
{21'b000000000000011100111, 21'b111111111110011001101, 21'b111111111110100011010, 21'b111111111111101010001, 21'b000000000001010101101, 21'b111111111111111111111, 21'b111111111111010011101, 21'b000000000000100001111, 21'b000000000000000111100, 21'b000000000000000000000, 21'b000000000000011010101, 21'b111111111111011101010, 21'b000000000000000000000, 21'b000000000000000000100, 21'b111111111111111011111, 21'b000000000000000010010, 21'b111111111111110010101, 21'b111111111110001010000, 21'b000000000000010101011, 21'b000000000000101100001, 21'b000000000000100001111, 21'b000000000000000000010, 21'b000000000000000011101, 21'b111111111111001100011, 21'b111111111110101111000, 21'b111111111111111111010, 21'b111111111111011001101, 21'b111111111111000101011, 21'b111111111111100111000, 21'b111111111110001111101, 21'b000000000000110101101, 21'b000000000000110110111}, 
{21'b000000000000000000000, 21'b000000000000000000000, 21'b000000000000000000010, 21'b000000000000000000000, 21'b000000000000100001001, 21'b111111111111101000000, 21'b000000000000000010010, 21'b000000000000001001010, 21'b111111111111010011010, 21'b000000000000000100101, 21'b111111111111111111011, 21'b111111111111111111111, 21'b111111111111111111111, 21'b000000000000011110101, 21'b000000000000000110101, 21'b000000000000000010110, 21'b000000000000000111111, 21'b000000000000101010101, 21'b111111111111100100000, 21'b000000000000000000000, 21'b111111111111101010111, 21'b111111111111111111111, 21'b000000000000101000010, 21'b000000000000000001000, 21'b111111111111111111101, 21'b111111111110111000001, 21'b111111111111111110110, 21'b111111111111101100001, 21'b111111111111111000001, 21'b000000000000000000011, 21'b000000000000010001010, 21'b000000000000001101010}, 
{21'b111111111111111010011, 21'b000000000000010001001, 21'b111111111111011001000, 21'b000000000000000010101, 21'b000000000000011000110, 21'b111111111111111010111, 21'b111111111111111111011, 21'b000000000000010100111, 21'b000000000000000000000, 21'b111111111111111111111, 21'b111111111111110111101, 21'b000000000000000000000, 21'b000000000000000000000, 21'b111111111111111011100, 21'b111111111111110000011, 21'b111111111111110111100, 21'b111111111111111000110, 21'b111111111111110111111, 21'b111111111111110001111, 21'b000000000000000000000, 21'b111111111111111111111, 21'b111111111111111010010, 21'b111111111111110111011, 21'b000000000000110010111, 21'b000000000000000000000, 21'b111111111111010001111, 21'b111111111111111110111, 21'b000000000000001111110, 21'b000000000000000000000, 21'b000000000000000000000, 21'b000000000000100000000, 21'b111111111111111111111}, 
{21'b111111111111111111111, 21'b000000000000000000100, 21'b111111111111111111111, 21'b111111111111101100000, 21'b111111111110010001111, 21'b000000000000000000000, 21'b000000000000000000000, 21'b111111111111111111001, 21'b111111111110110011010, 21'b000000000000001010011, 21'b111111111111110011011, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111010000101, 21'b111111111111111010001, 21'b111111111111111111111, 21'b000000000000000000001, 21'b000000000000000001000, 21'b000000000000000100101, 21'b000000000000101100001, 21'b111111111111110000101, 21'b111111111111011001101, 21'b000000000000000000000, 21'b111111111111011110111, 21'b111111111111110011010, 21'b111111111111100010011, 21'b111111111111111111000, 21'b111111111111111110011, 21'b111111111111111101101, 21'b111111111111000011101, 21'b111111111111111011101, 21'b000000000000011111000}, 
{21'b000000000000001110011, 21'b000000000000011100000, 21'b111111111111111111101, 21'b000000000000010100011, 21'b111111111111100101000, 21'b111111111111110000000, 21'b000000000000001100001, 21'b000000000000001000110, 21'b111111111111111001111, 21'b111111111111111111111, 21'b111111111111111111111, 21'b111111111111111111111, 21'b111111111111111111111, 21'b111111111111010110111, 21'b111111111111111111111, 21'b000000000000010010011, 21'b111111111111110001010, 21'b000000000000000100011, 21'b111111111111111111110, 21'b111111111111111111110, 21'b000000000000011010100, 21'b111111111111010110001, 21'b000000000000100011111, 21'b000000000000000110000, 21'b000000000000000000000, 21'b000000000000011011000, 21'b000000000000000000011, 21'b111111111111111011011, 21'b111111111111001111010, 21'b111111111111110001111, 21'b111111111111101010001, 21'b000000000000010110101}, 
{21'b000000000000000000000, 21'b000000000000000000111, 21'b111111111111010001001, 21'b111111111111111111101, 21'b000000000000011010011, 21'b111111111111101101111, 21'b111111111111111110011, 21'b111111111111111111111, 21'b000000000000000010100, 21'b000000000000000000000, 21'b000000000000000000000, 21'b111111111111100101111, 21'b000000000000001100010, 21'b000000000000000000110, 21'b000000000000000000000, 21'b000000000000000100110, 21'b111111111111111111111, 21'b111111111111101100111, 21'b000000000000000010010, 21'b000000000000000000000, 21'b111111111111111011100, 21'b111111111111111101001, 21'b000000000000100101111, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111011010100, 21'b111111111111010110001, 21'b000000000000011110111, 21'b111111111111111111110, 21'b111111111111111111111, 21'b000000000000000011100, 21'b000000000000100100001}, 
{21'b111111111111010100011, 21'b111111111111111111111, 21'b111111111111100100110, 21'b000000000000000000100, 21'b111111111111010010110, 21'b000000000000000000000, 21'b111111111111111111111, 21'b111111111111110111101, 21'b111111111110111011110, 21'b111111111111111100101, 21'b000000000000000000000, 21'b111111111111111110111, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111111110111, 21'b111111111111111001101, 21'b111111111111101101000, 21'b111111111111110011110, 21'b000000000000001000011, 21'b111111111111111111101, 21'b111111111111111100110, 21'b000000000000000000000, 21'b000000000000101011000, 21'b111111111111111111111, 21'b000000000000010011001, 21'b000000000000001011101, 21'b111111111111101110011, 21'b000000000000011011010, 21'b111111111111111010001, 21'b000000000000000000000, 21'b111111111111111111110, 21'b000000000001001010100}, 
{21'b111111111111010111110, 21'b000000000000000011110, 21'b000000000000000110011, 21'b111111111111111100011, 21'b000000000000011111010, 21'b111111111111011001010, 21'b111111111111111111000, 21'b000000000000100001111, 21'b000000000000010100011, 21'b000000000000000001001, 21'b111111111111111111111, 21'b111111111111110111001, 21'b111111111111110100100, 21'b111111111111110111101, 21'b111111111111111001101, 21'b000000000000001011100, 21'b111111111111111111111, 21'b000000000000000001000, 21'b000000000000010010000, 21'b000000000000000000000, 21'b000000000000000000000, 21'b000000000000000001111, 21'b000000000000100000010, 21'b000000000000000101110, 21'b000000000000000000110, 21'b111111111111110010001, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111111110001, 21'b111111111111111110011, 21'b111111111111111111111, 21'b000000000000001000101}, 
{21'b111111111111111111111, 21'b000000000000000000011, 21'b111111111111100100110, 21'b111111111111110110011, 21'b000000000000100100000, 21'b111111111111111111111, 21'b111111111111110110000, 21'b000000000000011111010, 21'b111111111111111001001, 21'b000000000000100101010, 21'b000000000000001010111, 21'b111111111111110000100, 21'b000000000000000000000, 21'b000000000000000000011, 21'b111111111111111110000, 21'b000000000000000010101, 21'b111111111111110110001, 21'b111111111111011110010, 21'b000000000000100011100, 21'b000000000000010011111, 21'b000000000001010001001, 21'b000000000000011001101, 21'b000000000000011111110, 21'b111111111111111111111, 21'b000000000000000000000, 21'b000000000000000000000, 21'b000000000000000111010, 21'b000000000000001010001, 21'b111111111111001010001, 21'b111111111111111111111, 21'b111111111111111111010, 21'b111111111111111111001}, 
{21'b000000000000000000000, 21'b111111111111110100110, 21'b111111111111110010101, 21'b000000000000000000000, 21'b111111111111100000110, 21'b000000000000000000000, 21'b000000000000011000100, 21'b000000000000001101111, 21'b000000000000000110110, 21'b111111111111110011010, 21'b000000000000000000000, 21'b111111111111111111111, 21'b111111111111111111111, 21'b111111111111111111111, 21'b111111111111111010100, 21'b000000000000011001110, 21'b111111111111111111111, 21'b111111111111111111111, 21'b111111111111011001010, 21'b000000000000000000000, 21'b111111111111100111010, 21'b111111111111111111110, 21'b000000000000000000000, 21'b111111111111111111011, 21'b000000000000000001111, 21'b000000000000000010001, 21'b000000000000000011100, 21'b000000000000010001101, 21'b111111111111110111101, 21'b111111111111111111000, 21'b111111111111000110100, 21'b000000000000001010000}, 
{21'b000000000000111000100, 21'b111111111111111110111, 21'b000000000000001000011, 21'b111111111111110010100, 21'b111111111111110101000, 21'b000000000000000100010, 21'b000000000000010100100, 21'b000000000000000000000, 21'b000000000001000011011, 21'b000000000000000000000, 21'b111111111111111101010, 21'b000000000000000010011, 21'b000000000000001100000, 21'b111111111111111111101, 21'b000000000000000110110, 21'b000000000000001101001, 21'b111111111111111111011, 21'b111111111111000111000, 21'b111111111111111000110, 21'b111111111111111111110, 21'b000000000000001110111, 21'b000000000000000000001, 21'b111111111111111111111, 21'b000000000000001110011, 21'b000000000000000010010, 21'b111111111111011110010, 21'b111111111111110010110, 21'b000000000000010000111, 21'b111111111111111100011, 21'b000000000000100001000, 21'b111111111111111111110, 21'b111111111111101001000}, 
{21'b000000000000000001101, 21'b000000000000001101000, 21'b111111111111111111111, 21'b111111111111111011000, 21'b111111111111010010110, 21'b111111111111111111111, 21'b000000000000000101111, 21'b111111111111111010000, 21'b000000000000010101000, 21'b111111111111111011101, 21'b111111111111111111111, 21'b111111111111111011101, 21'b111111111111111111111, 21'b111111111111111011010, 21'b000000000000000000000, 21'b000000000000101000000, 21'b000000000000000000000, 21'b111111111111111111110, 21'b111111111111111111111, 21'b111111111111111111111, 21'b111111111111111111111, 21'b111111111111111111111, 21'b000000000000000100010, 21'b000000000000010000000, 21'b000000000000000000000, 21'b000000000000000000100, 21'b000000000000000100001, 21'b111111111111111111111, 21'b000000000000000000000, 21'b000000000000000010100, 21'b000000000000000000001, 21'b000000000000001100011}, 
{21'b111111111111011000011, 21'b000000000000010000101, 21'b000000000000000010010, 21'b111111111111110010100, 21'b111111111111001100111, 21'b111111111111111101101, 21'b000000000000001000100, 21'b111111111111001101001, 21'b000000000001000001011, 21'b000000000000001001001, 21'b000000000000000010000, 21'b000000000000001100000, 21'b000000000000000101101, 21'b000000000000000000000, 21'b000000000000110100001, 21'b111111111111110101001, 21'b000000000000000000101, 21'b000000000000000000000, 21'b111111111111111111001, 21'b000000000000000000011, 21'b111111111111001000101, 21'b000000000000000010001, 21'b000000000000010011100, 21'b000000000000000100110, 21'b000000000000000100100, 21'b111111111110101011111, 21'b111111111111010100010, 21'b111111111111100001001, 21'b000000000000000000010, 21'b111111111111111111110, 21'b000000000000101001101, 21'b111111111111100101110}, 
{21'b111111111111111110010, 21'b111111111111100111000, 21'b111111111111110010110, 21'b111111111111001011101, 21'b111111111111011110101, 21'b000000000000101011000, 21'b000000000000100111101, 21'b111111111111101010001, 21'b000000000000000101010, 21'b111111111111111011000, 21'b111111111111110011111, 21'b111111111111011111110, 21'b000000000000001101001, 21'b111111111111011011101, 21'b000000000000011000001, 21'b111111111111111111111, 21'b000000000000101010111, 21'b111111111111111111111, 21'b111111111111111111000, 21'b111111111111101110101, 21'b111111111111111010101, 21'b111111111111110111101, 21'b111111111111011101111, 21'b000000000000001010100, 21'b111111111111111111111, 21'b111111111111111111001, 21'b111111111111100010110, 21'b000000000000101000010, 21'b000000000000100011101, 21'b111111111111110100011, 21'b111111111110101111010, 21'b000000000000010010010}, 
{21'b000000000000000000000, 21'b111111111111111100101, 21'b111111111111111111111, 21'b111111111111110011100, 21'b000000000000000011101, 21'b000000000000000001001, 21'b000000000000001000111, 21'b000000000000000000101, 21'b000000000000001111000, 21'b111111111111111111111, 21'b000000000000000000000, 21'b000000000000001100001, 21'b000000000000000000001, 21'b000000000000000001100, 21'b111111111111101111000, 21'b111111111111110010001, 21'b000000000000000000000, 21'b000000000000010111010, 21'b000000000000000111010, 21'b000000000000010000000, 21'b111111111111111101111, 21'b111111111111101011100, 21'b111111111111111111111, 21'b000000000000001001100, 21'b111111111111111111111, 21'b000000000000000100001, 21'b111111111111111111011, 21'b000000000000001000101, 21'b000000000000000000000, 21'b000000000000001010101, 21'b111111111111001111011, 21'b111111111111111111111}, 
{21'b000000000000100111101, 21'b111111111111111110110, 21'b000000000000010011001, 21'b111111111111011000111, 21'b111111111111100111010, 21'b111111111111111111111, 21'b111111111111111111111, 21'b000000000000000011100, 21'b000000000000000000010, 21'b111111111111101111111, 21'b000000000000000000000, 21'b000000000000000000010, 21'b000000000000000000000, 21'b000000000000000000000, 21'b111111111111101111011, 21'b000000000000010010010, 21'b111111111111111111110, 21'b111111111111111100000, 21'b000000000000000000000, 21'b000000000000001111010, 21'b111111111111100110010, 21'b000000000000001110110, 21'b000000000000010001111, 21'b000000000000010000100, 21'b111111111111111111111, 21'b000000000001000110100, 21'b111111111111101100011, 21'b000000000000101110100, 21'b111111111111111001011, 21'b111111111111010001110, 21'b111111111111101001110, 21'b000000000000010001110}, 
{21'b111111111110111010011, 21'b111111111111111100100, 21'b111111111111101100010, 21'b111111111111111111111, 21'b000000000000100001011, 21'b111111111111101001001, 21'b111111111111111000010, 21'b000000000000011110011, 21'b000000000000001100000, 21'b111111111111100001100, 21'b000000000000000000000, 21'b111111111111111100011, 21'b111111111111111110101, 21'b000000000000010001100, 21'b111111111111100000100, 21'b111111111111111110100, 21'b000000000000000000000, 21'b111111111111111111111, 21'b111111111111111101111, 21'b000000000000000000000, 21'b111111111111100111101, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111010101111, 21'b000000000000001000111, 21'b000000000001001111010, 21'b000000000000101100010, 21'b111111111111111011011, 21'b111111111111101011011, 21'b111111111111000110100, 21'b000000000000000000000, 21'b111111111111111001110}, 
{21'b000000000000000010101, 21'b000000000000011011010, 21'b000000000000000010101, 21'b111111111111101100101, 21'b000000000000000000100, 21'b111111111111111100101, 21'b000000000000000000000, 21'b000000000000011010101, 21'b000000000000011011100, 21'b111111111111101110111, 21'b000000000000010001111, 21'b000000000000000011000, 21'b111111111111111111111, 21'b111111111111111110001, 21'b111111111111101011101, 21'b000000000000100000011, 21'b111111111111111010100, 21'b111111111111010110101, 21'b000000000000001110101, 21'b111111111111111111111, 21'b111111111111111111111, 21'b000000000000001110111, 21'b111111111111110110011, 21'b111111111111111111011, 21'b111111111111111001011, 21'b000000000000001011010, 21'b111111111111101110000, 21'b000000000000010001001, 21'b111111111111010001011, 21'b000000000000001010010, 21'b111111111111111111111, 21'b000000000000010100000}, 
{21'b111111111111111010100, 21'b000000000000000000000, 21'b000000000000001011011, 21'b000000000000000000000, 21'b111111111111111000001, 21'b111111111111111111101, 21'b000000000000001101001, 21'b111111111111111111111, 21'b000000000000000000000, 21'b000000000000000000101, 21'b000000000000000000000, 21'b000000000000000010100, 21'b111111111111110010011, 21'b000000000000000001010, 21'b000000000000001110001, 21'b000000000000000101111, 21'b000000000000001101100, 21'b111111111111111111111, 21'b111111111111111111110, 21'b000000000000010000011, 21'b000000000000011111101, 21'b111111111111110011011, 21'b000000000000000000000, 21'b111111111111111111101, 21'b000000000000000001011, 21'b111111111111000100111, 21'b111111111111111111111, 21'b111111111111110110111, 21'b111111111111111111111, 21'b000000000001001000010, 21'b000000000000000000000, 21'b111111111111100101101}, 
{21'b111111111111111100100, 21'b111111111111110000101, 21'b111111111111111110110, 21'b000000000000000000111, 21'b000000000000001011100, 21'b111111111111111111111, 21'b000000000000000000000, 21'b111111111111111101000, 21'b000000000000001001000, 21'b111111111111111110111, 21'b000000000000000000000, 21'b000000000000000100000, 21'b000000000000100101110, 21'b111111111111110010111, 21'b000000000000000001100, 21'b111111111110010011011, 21'b111111111111111110100, 21'b111111111111111000010, 21'b000000000000000001000, 21'b111111111111111001100, 21'b000000000000001011110, 21'b111111111111100011010, 21'b000000000000001110100, 21'b000000000000001101011, 21'b111111111111111110010, 21'b111111111110100100111, 21'b111111111111100010101, 21'b111111111111111101001, 21'b111111111111111101101, 21'b000000000000110001111, 21'b111111111111111111010, 21'b000000000000010011101}, 
{21'b000000000000000110000, 21'b000000000000000000000, 21'b000000000000010110010, 21'b111111111111110001011, 21'b111111111111110111001, 21'b000000000000011110011, 21'b111111111111101011100, 21'b000000000000000111010, 21'b111111111111011000011, 21'b000000000000000001000, 21'b000000000000000010001, 21'b111111111111110101010, 21'b000000000000000000000, 21'b000000000000000000000, 21'b111111111111100111111, 21'b000000000000110111010, 21'b111111111111100000011, 21'b111111111111111110011, 21'b000000000000001111001, 21'b111111111111111111111, 21'b000000000000001000110, 21'b111111111111000010101, 21'b000000000000101000000, 21'b111111111111111111111, 21'b111111111111110000001, 21'b000000000000111110000, 21'b000000000000010010101, 21'b111111111111101011110, 21'b111111111111101110110, 21'b111111111110111011001, 21'b111111111111111110101, 21'b000000000000000010000}, 
{21'b111111111111111111111, 21'b000000000000000000110, 21'b111111111111111011100, 21'b111111111111011101101, 21'b111111111111111111111, 21'b111111111111001101110, 21'b000000000000000000000, 21'b000000000000100110110, 21'b000000000000011111010, 21'b000000000000000010011, 21'b000000000000000000000, 21'b111111111111110001111, 21'b000000000000101010100, 21'b111111111111111111111, 21'b111111111111111111111, 21'b111111111111111111111, 21'b000000000000110111100, 21'b000000000000000000001, 21'b111111111111111010111, 21'b111111111111111001011, 21'b111111111111010110110, 21'b000000000000010000110, 21'b000000000000000000000, 21'b000000000000000000000, 21'b000000000000000100000, 21'b111111111111110110111, 21'b111111111111000101000, 21'b000000000000100011010, 21'b111111111111000111001, 21'b000000000000000110100, 21'b111111111111110101111, 21'b000000000000000000000}, 
{21'b000000000000000111110, 21'b000000000000010111110, 21'b000000000000000001001, 21'b111111111111111111100, 21'b111111111111000101001, 21'b000000000000000000000, 21'b111111111111111111111, 21'b000000000000011111000, 21'b000000000000100011011, 21'b111111111111111111111, 21'b111111111111111111111, 21'b111111111111111111110, 21'b000000000000000000000, 21'b000000000000000000010, 21'b000000000000000000000, 21'b000000000000000000000, 21'b000000000000000000000, 21'b111111111111111111111, 21'b000000000000010101110, 21'b111111111111110010110, 21'b111111111111001000101, 21'b111111111111111011110, 21'b111111111111110011010, 21'b111111111111110011111, 21'b111111111111110111001, 21'b111111111111111111111, 21'b111111111111110111111, 21'b111111111111111101001, 21'b111111111111111110101, 21'b000000000000010010000, 21'b111111111111111111111, 21'b000000000000111011010}
};

localparam logic signed [20:0] bias [32] = '{
21'b000000000010111100101,  // 1.474280834197998
21'b000000000001011000100,  // 0.6914801001548767
21'b000000000010111000011,  // 1.4406442642211914
21'b000000000010110100001,  // 1.408045768737793
21'b000000000001111110010,  // 0.9864811301231384
21'b000000000001101110100,  // 0.8636202812194824
21'b111111111110110001001,  // -0.6153604388237
21'b000000000000111101111,  // 0.4839226007461548
21'b000000000000111110001,  // 0.4862793982028961
21'b000000000000101111100,  // 0.37162142992019653
21'b000000000000111010110,  // 0.45989668369293213
21'b000000000010100110011,  // 1.2998151779174805
21'b111111111101111101111,  // -1.016528844833374
21'b111111111111010010111,  // -0.35249894857406616
21'b000000000000111001000,  // 0.44582197070121765
21'b111111111111110001101,  // -0.1119980737566948
21'b111111111111110111011,  // -0.06717441976070404
21'b000000000000000000100,  // 0.00487547367811203
21'b000000000000011000111,  // 0.1946917623281479
21'b111111111110011100001,  // -0.7796769738197327
21'b000000000001011101010,  // 0.7287401556968689
21'b000000000011011011100,  // 1.714877724647522
21'b111111111100110011100,  // -1.5971007347106934
21'b000000000000001001011,  // 0.07393483817577362
21'b000000000000101001010,  // 0.3225609362125397
21'b000000000001101100001,  // 0.8453295230865479
21'b000000000001110011000,  // 0.898597240447998
21'b000000000000100000100,  // 0.2548799514770508
21'b000000000001111100100,  // 0.9735668301582336
21'b000000000010010000001,  // 1.1261906623840332
21'b000000000000111001010,  // 0.44768181443214417
21'b111111111011010000111   // -2.3676068782806396
};
endpackage