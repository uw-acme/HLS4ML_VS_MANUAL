// Width: 15
// NFRAC: 7
package dense_2_15_7;

localparam logic signed [14:0] weights [64][32] = '{ 
{15'b000000000100010, 15'b000000000000001, 15'b111111111100111, 15'b111111111111101, 15'b000000000100001, 15'b000000000000000, 15'b111111111101101, 15'b111111111111111, 15'b111111111011100, 15'b000000000001010, 15'b000000000000000, 15'b111111111111111, 15'b111111111111111, 15'b111111111100110, 15'b111111111111001, 15'b111111111011110, 15'b000000000000000, 15'b111111111111110, 15'b111111111100111, 15'b111111111101011, 15'b000000000000000, 15'b000000000000000, 15'b111111111111110, 15'b111111111111111, 15'b000000000000000, 15'b000000000001100, 15'b000000000110001, 15'b000000000010110, 15'b111111111111111, 15'b000000000000110, 15'b111111111001011, 15'b000000000000000}, 
{15'b111111111110011, 15'b111111111101100, 15'b111111111101110, 15'b111111111111000, 15'b111111111111111, 15'b000000000000101, 15'b111111111100011, 15'b000000000000000, 15'b000000000000000, 15'b111111111110111, 15'b000000000010011, 15'b111111111111010, 15'b111111111111000, 15'b111111111100100, 15'b000000000000000, 15'b111111111111001, 15'b000000000000001, 15'b111111111100111, 15'b000000000010101, 15'b000000000011101, 15'b111111111111011, 15'b111111111111111, 15'b111111111111111, 15'b000000000000011, 15'b111111111110110, 15'b000000000100011, 15'b000000000011111, 15'b000000000000001, 15'b000000000000011, 15'b111111111000001, 15'b000000000000000, 15'b000000000000000}, 
{15'b000000000001001, 15'b111111111110001, 15'b111111111101111, 15'b111111111111010, 15'b111111111110110, 15'b111111111110101, 15'b111111111101000, 15'b000000000000000, 15'b111111111101110, 15'b000000000000001, 15'b000000000000000, 15'b111111111110101, 15'b000000000001011, 15'b111111111110111, 15'b111111111111111, 15'b111111111111011, 15'b000000000000000, 15'b000000000001100, 15'b000000000000111, 15'b000000000011101, 15'b000000000000101, 15'b111111111110101, 15'b000000000000000, 15'b000000000000100, 15'b111111111111101, 15'b000000000011010, 15'b000000000010011, 15'b000000000001100, 15'b111111111111111, 15'b111111111101100, 15'b111111111111110, 15'b000000000001100}, 
{15'b000000000010001, 15'b000000000000010, 15'b000000000000110, 15'b111111111111110, 15'b111111110111110, 15'b000000000000000, 15'b000000000000000, 15'b000000000011100, 15'b000000000011111, 15'b111111111111110, 15'b111111111111111, 15'b000000000000000, 15'b000000000000000, 15'b000000000000000, 15'b111111111111101, 15'b000000000011011, 15'b000000000000000, 15'b111111111111100, 15'b111111111111111, 15'b111111111101001, 15'b111111111111000, 15'b000000000000110, 15'b111111111110111, 15'b111111111111111, 15'b000000000000000, 15'b111111111111001, 15'b000000000001001, 15'b111111111111111, 15'b111111111111111, 15'b111111111111111, 15'b111111111100100, 15'b000000000100111}, 
{15'b111111110101000, 15'b111111111111100, 15'b111111111111111, 15'b000000000000000, 15'b111111111111100, 15'b000000000000000, 15'b111111111111001, 15'b111111111101100, 15'b000000000000110, 15'b111111111111101, 15'b111111111111110, 15'b111111111111111, 15'b111111111111111, 15'b000000000011010, 15'b000000000000000, 15'b000000000101010, 15'b111111111111111, 15'b000000000011011, 15'b111111111001100, 15'b000000000000000, 15'b111111111110001, 15'b000000000010101, 15'b000000000100001, 15'b000000000000000, 15'b000000000000101, 15'b000000000010100, 15'b000000000011110, 15'b000000000000010, 15'b111111111111111, 15'b111111111111111, 15'b111111111111110, 15'b000000000011100}, 
{15'b000000000000111, 15'b111111111111111, 15'b000000000010011, 15'b111111110101100, 15'b111111101001111, 15'b111111111010011, 15'b000000000101101, 15'b111111110110000, 15'b111111111111111, 15'b111111110101001, 15'b111111110111111, 15'b111111111010100, 15'b000000000101101, 15'b111111111111111, 15'b111111111111110, 15'b000000000000000, 15'b111111111111111, 15'b111111111111111, 15'b111111111101111, 15'b111111111111111, 15'b111111111000001, 15'b000000000000000, 15'b000000000010111, 15'b111111111111111, 15'b000000000000010, 15'b000000000100010, 15'b000000000000110, 15'b111111111111111, 15'b111111111111111, 15'b000000000011010, 15'b111111111111011, 15'b000000000011001}, 
{15'b111111111111011, 15'b111111111101011, 15'b111111111100001, 15'b111111111111001, 15'b111111111011011, 15'b000000000001000, 15'b111111111101000, 15'b111111111101101, 15'b111111111001010, 15'b000000000000110, 15'b111111111111111, 15'b111111111101011, 15'b000000000001111, 15'b111111111111110, 15'b111111111111010, 15'b111111110111001, 15'b111111111111111, 15'b000000000001010, 15'b000000000011000, 15'b111111111101011, 15'b111111111101100, 15'b111111111110111, 15'b111111111111111, 15'b000000000000011, 15'b111111111111010, 15'b111111110101101, 15'b111111111011110, 15'b111111111111010, 15'b000000000000000, 15'b111111111111101, 15'b000000000000011, 15'b111111111111111}, 
{15'b111111111101100, 15'b111111111110100, 15'b111111111110101, 15'b111111111100001, 15'b111111111110001, 15'b111111111111111, 15'b000000000001101, 15'b111111111110101, 15'b000000000011001, 15'b000000000000000, 15'b000000000000000, 15'b111111111111111, 15'b000000000011100, 15'b000000000000000, 15'b111111111111111, 15'b111111111110110, 15'b111111111111111, 15'b000000000000000, 15'b111111111111111, 15'b000000000000000, 15'b111111111111111, 15'b111111111111111, 15'b000000000000000, 15'b111111111111111, 15'b000000000000101, 15'b111111111101000, 15'b000000000000001, 15'b111111111111111, 15'b111111111110110, 15'b111111111111111, 15'b000000000000000, 15'b111111111111111}, 
{15'b111111111000010, 15'b111111111111000, 15'b111111111001111, 15'b000000000001111, 15'b000000000111110, 15'b111111111111111, 15'b111111111111100, 15'b000000000011110, 15'b111111111000111, 15'b111111111111010, 15'b000000000000000, 15'b111111111100110, 15'b111111111111111, 15'b000000000001001, 15'b111111111100111, 15'b000000001100000, 15'b111111111111110, 15'b000000000000101, 15'b000000000011010, 15'b000000000011111, 15'b000000000000000, 15'b111111111010101, 15'b000000000000000, 15'b000000000110100, 15'b111111111101000, 15'b000000001011001, 15'b111111111101100, 15'b111111111100101, 15'b111111111000011, 15'b111111111000100, 15'b000000000000000, 15'b000000000000110}, 
{15'b000000000000000, 15'b111111111111110, 15'b111111111110110, 15'b000000000000000, 15'b000000000100111, 15'b111111111111101, 15'b111111111110111, 15'b000000000001011, 15'b000000000001100, 15'b000000000000000, 15'b111111111111110, 15'b111111111111111, 15'b111111111111111, 15'b111111111110001, 15'b111111111111111, 15'b000000000000000, 15'b000000000000000, 15'b111111111111111, 15'b000000000000000, 15'b000000000001010, 15'b000000000000010, 15'b111111111111111, 15'b000000000000000, 15'b000000000000000, 15'b000000000000100, 15'b111111111101111, 15'b000000000001000, 15'b000000000011111, 15'b111111111111111, 15'b000000000000000, 15'b000000000000110, 15'b000000000001000}, 
{15'b000000000001100, 15'b000000000000000, 15'b111111111110010, 15'b111111111011111, 15'b111111110011010, 15'b000000000010001, 15'b000000000000000, 15'b111111110010110, 15'b000000000000100, 15'b111111111111111, 15'b000000000000000, 15'b111111111111111, 15'b000000000000001, 15'b000000000000000, 15'b111111111111101, 15'b111111111001111, 15'b111111111111111, 15'b000000000011100, 15'b000000000010000, 15'b000000000011000, 15'b111111111000111, 15'b111111111010010, 15'b000000000001111, 15'b111111111111011, 15'b111111111111010, 15'b000000000101101, 15'b111111111110011, 15'b111111111111111, 15'b111111111111111, 15'b000000000011011, 15'b111111111111111, 15'b000000000000000}, 
{15'b111111111100110, 15'b111111111000000, 15'b000000000000000, 15'b111111111111111, 15'b000000000101010, 15'b111111111011101, 15'b111111111100011, 15'b000000000001110, 15'b111111111111111, 15'b000000000010011, 15'b000000000001001, 15'b111111111110110, 15'b000000000000000, 15'b000000000000001, 15'b111111111111101, 15'b111111111011111, 15'b000000000010110, 15'b000000000000011, 15'b000000000100110, 15'b000000000001011, 15'b000000000000000, 15'b111111111111011, 15'b000000000010000, 15'b111111111110100, 15'b111111111011000, 15'b111111111111111, 15'b000000000010111, 15'b111111111111111, 15'b000000000000001, 15'b111111111110011, 15'b000000000010001, 15'b000000000100011}, 
{15'b000000000000001, 15'b000000000000000, 15'b000000000011100, 15'b000000000000001, 15'b111111111111010, 15'b000000000010111, 15'b000000000001011, 15'b111111111111111, 15'b000000000000000, 15'b111111111101110, 15'b111111111111001, 15'b111111111101010, 15'b111111111111111, 15'b000000000000110, 15'b111111111110111, 15'b000000001101011, 15'b000000000000000, 15'b111111111110011, 15'b111111111100111, 15'b111111111111110, 15'b000000000011001, 15'b000000000010000, 15'b000000000000000, 15'b111111111111111, 15'b000000000011100, 15'b000000000100010, 15'b000000000111111, 15'b000000000000001, 15'b000000000000000, 15'b000000000000000, 15'b111111111111110, 15'b111111111110110}, 
{15'b111111111101100, 15'b000000000000110, 15'b000000000000101, 15'b111111111100000, 15'b111111111011101, 15'b000000000111100, 15'b000000000000110, 15'b000000000000000, 15'b111111111101011, 15'b111111111110100, 15'b000000000010000, 15'b000000000001001, 15'b000000000000000, 15'b111111111110101, 15'b000000000100100, 15'b111111111111111, 15'b111111111111110, 15'b000000000000000, 15'b000000000000001, 15'b111111111111010, 15'b000000000001010, 15'b000000000000010, 15'b000000000001110, 15'b111111111111111, 15'b000000000000000, 15'b000000001010100, 15'b111111111111000, 15'b111111111111101, 15'b111111111111111, 15'b111111111110010, 15'b111111111111010, 15'b000000000010110}, 
{15'b000000000000111, 15'b000000000001001, 15'b000000000101001, 15'b111111111111010, 15'b000000000001100, 15'b000000000101100, 15'b000000000000000, 15'b111111111111100, 15'b000000000001111, 15'b111111111110001, 15'b111111111111111, 15'b111111111110000, 15'b000000000000000, 15'b000000000110010, 15'b111111111111101, 15'b000000000000000, 15'b000000000011110, 15'b000000000000000, 15'b000000000000000, 15'b111111111010111, 15'b111111111100000, 15'b111111111111011, 15'b111111111111111, 15'b111111111101101, 15'b111111111111011, 15'b111111111110101, 15'b111111111100110, 15'b111111111100100, 15'b000000000000011, 15'b000000000001110, 15'b111111111001101, 15'b000000000000000}, 
{15'b111111111011001, 15'b000000000000000, 15'b111111111111110, 15'b111111111111001, 15'b111111111111111, 15'b000000000010001, 15'b111111111110110, 15'b000000000100010, 15'b111111111010001, 15'b111111111111111, 15'b000000000000000, 15'b111111111111111, 15'b000000000000000, 15'b000000000000000, 15'b111111111111111, 15'b111111111110100, 15'b000000000001010, 15'b000000000010111, 15'b111111111111110, 15'b111111111011111, 15'b111111111111000, 15'b000000000001110, 15'b000000000001000, 15'b000000000000000, 15'b000000000000000, 15'b000000000001010, 15'b111111111100001, 15'b000000000000000, 15'b111111111111111, 15'b000000000000000, 15'b000000000000000, 15'b111111111101111}, 
{15'b111111111010100, 15'b111111111111111, 15'b111111111111111, 15'b111111111111101, 15'b111111111111111, 15'b000000000001101, 15'b000000000000000, 15'b000000000000100, 15'b000000000000100, 15'b000000000001000, 15'b000000000001010, 15'b000000000010100, 15'b000000000000011, 15'b111111111110011, 15'b000000000000000, 15'b000000000110000, 15'b000000000000000, 15'b000000000000000, 15'b111111111111111, 15'b000000000001110, 15'b000000000010010, 15'b000000000000011, 15'b000000000000101, 15'b111111111111100, 15'b111111111111011, 15'b000000000000011, 15'b111111111110111, 15'b111111111101111, 15'b000000000011010, 15'b111111111111100, 15'b000000000000100, 15'b111111111100111}, 
{15'b000000000000000, 15'b111111111111111, 15'b000000000000100, 15'b000000000000000, 15'b000000001110100, 15'b111111111111111, 15'b000000000000000, 15'b111111111111111, 15'b000000000001110, 15'b111111111110110, 15'b000000000000000, 15'b000000000000000, 15'b000000000000000, 15'b000000000010000, 15'b000000000000000, 15'b111111111101101, 15'b111111111111111, 15'b111111111110111, 15'b000000000101001, 15'b000000000000000, 15'b111111111111111, 15'b111111111111111, 15'b000000000000000, 15'b111111111111111, 15'b000000000000000, 15'b000000000001000, 15'b000000000000000, 15'b000000000000000, 15'b111111111111111, 15'b111111111111111, 15'b000000000000000, 15'b000000000000101}, 
{15'b111111111111111, 15'b000000000000011, 15'b111111111111111, 15'b000000000000110, 15'b111111111111010, 15'b111111111110000, 15'b111111111111000, 15'b000000000100011, 15'b000000000000000, 15'b000000000001100, 15'b111111111111110, 15'b000000000001000, 15'b111111111111011, 15'b111111111101011, 15'b111111111100111, 15'b000000000000001, 15'b111111111111111, 15'b111111111111011, 15'b000000000000000, 15'b000000000000000, 15'b111111111111111, 15'b000000000001001, 15'b000000000000100, 15'b111111111101111, 15'b000000000001110, 15'b111111111101010, 15'b000000000000000, 15'b000000000000000, 15'b111111111101010, 15'b000000000000000, 15'b000000000000101, 15'b111111111111100}, 
{15'b111111111111110, 15'b111111111110011, 15'b000000000000000, 15'b111111111111000, 15'b000000000011011, 15'b111111111111111, 15'b111111111111101, 15'b000000000001101, 15'b111111111001101, 15'b000000000000000, 15'b111111111111011, 15'b111111111111111, 15'b000000000101100, 15'b000000000011101, 15'b111111111110011, 15'b111111111111101, 15'b111111111111111, 15'b000000000000000, 15'b111111111111111, 15'b000000000000000, 15'b000000000000000, 15'b111111111101110, 15'b111111111110000, 15'b000000000010000, 15'b000000000000000, 15'b111111111101110, 15'b000000000000011, 15'b111111111110101, 15'b111111111111011, 15'b000000000010001, 15'b000000000000000, 15'b111111111100000}, 
{15'b000000001010001, 15'b000000000101011, 15'b111111111100000, 15'b000000000000000, 15'b111111111010011, 15'b000000000000000, 15'b000000000011100, 15'b000000000000011, 15'b000000000011100, 15'b111111111111111, 15'b111111111101100, 15'b111111111110101, 15'b000000000010010, 15'b000000000000011, 15'b111111111110011, 15'b000000000010000, 15'b000000001000100, 15'b111111111101111, 15'b111111111011010, 15'b000000000000000, 15'b111111111111100, 15'b111111111101001, 15'b111111111111110, 15'b111111111111111, 15'b000000000001011, 15'b111111111010001, 15'b000000000001011, 15'b111111111111111, 15'b000000000000000, 15'b000000000001101, 15'b111111111111100, 15'b000000000000111}, 
{15'b111111111110100, 15'b111111111100111, 15'b111111111111011, 15'b111111111101010, 15'b111111111111101, 15'b000000000000110, 15'b000000000000000, 15'b111111111111110, 15'b000000000000100, 15'b111111111111111, 15'b000000000000000, 15'b111111111100100, 15'b000000000001101, 15'b000000000001010, 15'b111111111110010, 15'b000000000111000, 15'b111111111111111, 15'b000000000000000, 15'b111111111111111, 15'b000000000000000, 15'b000000000101000, 15'b111111111000011, 15'b111111111110010, 15'b111111111111000, 15'b111111111111101, 15'b000000000011001, 15'b111111111111001, 15'b000000000000010, 15'b000000000111101, 15'b111111110111110, 15'b111111111010001, 15'b000000000000010}, 
{15'b000000000000010, 15'b111111111111000, 15'b111111111111111, 15'b000000000000000, 15'b111111110100011, 15'b111111110110010, 15'b000000000000000, 15'b111111111111111, 15'b111111111011110, 15'b000000000000011, 15'b000000000000000, 15'b111111111111100, 15'b000000000000000, 15'b111111111111000, 15'b111111111111001, 15'b111111111110111, 15'b111111111101101, 15'b000000000100100, 15'b000000000000000, 15'b000000000000101, 15'b111111111111111, 15'b111111111110110, 15'b000000000000000, 15'b111111111110100, 15'b000000000011100, 15'b111111110110000, 15'b000000000011100, 15'b111111111111111, 15'b111111111111111, 15'b000000000011001, 15'b111111111111111, 15'b000000000011110}, 
{15'b111111111111111, 15'b000000000000000, 15'b111111111111010, 15'b000000000001001, 15'b000000000000111, 15'b111111111010100, 15'b000000000000000, 15'b000000000001000, 15'b000000001001010, 15'b111111111111110, 15'b000000000000000, 15'b000000000000111, 15'b000000000101101, 15'b111111111111011, 15'b000000000000001, 15'b000000000001100, 15'b111111111111111, 15'b000000000000011, 15'b111111111111111, 15'b000000000000000, 15'b111111111011100, 15'b000000000000100, 15'b000000000001000, 15'b000000000000010, 15'b111111111111111, 15'b000000000011011, 15'b000000000000000, 15'b000000000010000, 15'b111111111001010, 15'b000000000001101, 15'b000000000110010, 15'b000000000000000}, 
{15'b111111111010011, 15'b000000000011011, 15'b111111111011110, 15'b000000000001111, 15'b111111111110010, 15'b000000000000000, 15'b000000000111111, 15'b111111111100010, 15'b111111111011010, 15'b000000000010101, 15'b111111111100011, 15'b111111111111100, 15'b111111111111111, 15'b000000000101100, 15'b111111111111111, 15'b111111111011001, 15'b111111111111111, 15'b000000000111000, 15'b111111111000011, 15'b111111111111100, 15'b000000000101000, 15'b111111111010001, 15'b000000000000110, 15'b111111111111110, 15'b000000000100010, 15'b111111110111110, 15'b111111111010001, 15'b111111111100110, 15'b111111111111111, 15'b000000000001101, 15'b000000000000011, 15'b000000000010110}, 
{15'b111111111110100, 15'b000000000000110, 15'b111111111111111, 15'b000000000010011, 15'b111111111111011, 15'b000000000011101, 15'b000000000000000, 15'b111111111111110, 15'b111111111111111, 15'b000000000000000, 15'b000000000000000, 15'b111111111111111, 15'b111111111111111, 15'b000000001000010, 15'b000000000000001, 15'b000000000011000, 15'b000000000000000, 15'b111111111100100, 15'b111111111110110, 15'b111111111111111, 15'b111111111111101, 15'b000000000000101, 15'b111111111111111, 15'b111111111101000, 15'b111111111111111, 15'b000000000100101, 15'b000000000100111, 15'b111111111111111, 15'b111111111111101, 15'b000000000000000, 15'b111111111111111, 15'b111111111110011}, 
{15'b111111111110101, 15'b000000000000000, 15'b000000000100010, 15'b000000000000000, 15'b000000000000000, 15'b111111111110001, 15'b000000000000000, 15'b111111110010001, 15'b000000000011011, 15'b000000000000001, 15'b000000000000011, 15'b111111111010001, 15'b000000000000000, 15'b111111111101110, 15'b111111111111011, 15'b000000000000000, 15'b000000000000010, 15'b000000000000000, 15'b000000000001110, 15'b000000000000000, 15'b111111111111110, 15'b000000000101010, 15'b000000000110000, 15'b111111111100011, 15'b111111111101101, 15'b000000000011111, 15'b111111111011000, 15'b000000000000011, 15'b111111111111111, 15'b111111111111111, 15'b111111111111111, 15'b000000000010111}, 
{15'b111111111110001, 15'b111111111111111, 15'b111111111100001, 15'b111111111100110, 15'b111111111111110, 15'b111111111101110, 15'b000000000000000, 15'b000000000001011, 15'b111111111100001, 15'b111111111110101, 15'b111111111111001, 15'b000000000000000, 15'b000000000000011, 15'b111111111111110, 15'b111111111111000, 15'b000000000001100, 15'b000000000011100, 15'b000000000010000, 15'b111111111101111, 15'b000000000000110, 15'b111111111111110, 15'b111111111111100, 15'b000000000000010, 15'b000000000000010, 15'b111111111110111, 15'b000000000001011, 15'b111111111110100, 15'b000000000000111, 15'b111111111111111, 15'b111111111011010, 15'b111111111111100, 15'b000000000011100}, 
{15'b111111111111100, 15'b111111111110101, 15'b000000000001001, 15'b000000000100000, 15'b000000000001010, 15'b000000000001010, 15'b000000000000101, 15'b111111111100110, 15'b111111111100101, 15'b000000000001000, 15'b000000000000001, 15'b000000000000101, 15'b000000000000010, 15'b000000000000000, 15'b000000000011010, 15'b000000000000000, 15'b111111111111001, 15'b000000000001101, 15'b111111111111100, 15'b111111111111011, 15'b000000000001110, 15'b111111111110000, 15'b111111111111100, 15'b000000000010000, 15'b000000000000010, 15'b111111111110010, 15'b111111111100110, 15'b111111111111110, 15'b111111111011100, 15'b000000000000111, 15'b000000000001101, 15'b000000000000000}, 
{15'b111111111111110, 15'b111111111111101, 15'b111111111111110, 15'b111111111111011, 15'b111111111101111, 15'b111111111101110, 15'b000000000001000, 15'b000000000000001, 15'b111111111101000, 15'b000000000010101, 15'b111111111111101, 15'b111111111111111, 15'b111111111110001, 15'b000000000000000, 15'b000000000000011, 15'b111111111111001, 15'b111111111111101, 15'b111111111111010, 15'b111111111110101, 15'b000000000000000, 15'b111111111101110, 15'b000000000001101, 15'b111111111100100, 15'b000000000000000, 15'b000000000000101, 15'b000000000001111, 15'b000000000000011, 15'b000000000000000, 15'b000000000100101, 15'b000000000000110, 15'b000000000000000, 15'b000000000001010}, 
{15'b111111111111101, 15'b000000000100000, 15'b111111111111111, 15'b111111111111011, 15'b111111111100100, 15'b111111111110110, 15'b000000000110100, 15'b111111110100111, 15'b111111111010011, 15'b111111111100110, 15'b111111111100011, 15'b111111111011111, 15'b111111111111111, 15'b000000000111101, 15'b111111111111100, 15'b000000000000000, 15'b111111111100100, 15'b000000000111001, 15'b111111111001011, 15'b000000000000000, 15'b111111111111111, 15'b111111111010100, 15'b000000000000000, 15'b111111111111111, 15'b000000000000111, 15'b111111111111000, 15'b111111111101101, 15'b111111111111111, 15'b000000000010110, 15'b000000000000000, 15'b111111111110101, 15'b000000000000000}, 
{15'b000000000101111, 15'b111111111110001, 15'b000000000010000, 15'b111111111111011, 15'b000000000001001, 15'b111111111111111, 15'b111111111111111, 15'b111111111110100, 15'b000000000000000, 15'b000000000001011, 15'b111111111111111, 15'b111111111111000, 15'b111111111111111, 15'b000000000011101, 15'b000000000000010, 15'b000000000000101, 15'b000000000000011, 15'b111111111111100, 15'b000000000000010, 15'b000000000000000, 15'b111111111111110, 15'b111111111111111, 15'b111111111011000, 15'b111111111111111, 15'b000000000000111, 15'b111111111110001, 15'b111111111101110, 15'b111111111111111, 15'b111111111111111, 15'b000000001000111, 15'b111111111011011, 15'b111111111110001}, 
{15'b111111111111010, 15'b111111111110010, 15'b111111111110111, 15'b000000000000100, 15'b000000000010001, 15'b111111111101111, 15'b111111111111111, 15'b111111111100011, 15'b000000000000111, 15'b000000000010001, 15'b111111111100100, 15'b111111111011111, 15'b000000000000011, 15'b111111110101000, 15'b111111111110110, 15'b111111111110000, 15'b111111111100110, 15'b111111111111111, 15'b000000000010001, 15'b000000000000000, 15'b111111111111010, 15'b111111111111010, 15'b000000000000000, 15'b000000000000000, 15'b111111111111000, 15'b111111110011111, 15'b111111110111000, 15'b111111111011101, 15'b000000000000111, 15'b000000000011010, 15'b111111111111111, 15'b000000000011110}, 
{15'b111111111110100, 15'b111111111100100, 15'b000000000010100, 15'b000000000001001, 15'b000000000000101, 15'b111111111110100, 15'b111111111111011, 15'b000000000001100, 15'b000000001000100, 15'b111111111101010, 15'b111111111111111, 15'b111111111111111, 15'b000000000001111, 15'b111111111111000, 15'b111111111111101, 15'b111111111111101, 15'b111111111110011, 15'b111111111111111, 15'b000000000000000, 15'b000000000011101, 15'b111111111101110, 15'b111111111111111, 15'b000000000010000, 15'b111111111111110, 15'b000000000000000, 15'b000000001000011, 15'b000000000101001, 15'b000000000000000, 15'b000000000000000, 15'b111111111001010, 15'b111111111110111, 15'b111111111111111}, 
{15'b000000000000001, 15'b000000000000110, 15'b111111111111110, 15'b000000000000000, 15'b000000000011101, 15'b111111111000010, 15'b000000000000000, 15'b111111111110011, 15'b000000000010111, 15'b000000000000000, 15'b111111111111101, 15'b000000000000000, 15'b000000000000000, 15'b111111111111111, 15'b000000000000000, 15'b111111111110010, 15'b000000000100001, 15'b111111111111111, 15'b111111111111110, 15'b111111111111111, 15'b000000000000000, 15'b111111111111111, 15'b000000000000000, 15'b111111111111111, 15'b000000000000001, 15'b111111111010111, 15'b000000000000110, 15'b000000000010111, 15'b111111111111111, 15'b000000000001100, 15'b111111111111111, 15'b000000000001001}, 
{15'b111111111100110, 15'b000000000000001, 15'b111111111000010, 15'b000000000000000, 15'b111111111111001, 15'b111111111111010, 15'b111111111111111, 15'b111111111110100, 15'b111111111111011, 15'b111111111110111, 15'b000000000000110, 15'b000000000000011, 15'b111111111101001, 15'b000000000000000, 15'b111111111111111, 15'b111111111111110, 15'b000000000001001, 15'b111111111111101, 15'b111111111111100, 15'b111111111111100, 15'b111111111111111, 15'b000000000100010, 15'b111111111111111, 15'b000000000000000, 15'b111111111111110, 15'b000000000101000, 15'b000000000011000, 15'b000000000000100, 15'b111111111110011, 15'b111111111111110, 15'b000000000001000, 15'b000000000000111}, 
{15'b000000000000100, 15'b000000000000101, 15'b111111111111111, 15'b000000000000000, 15'b111111111000100, 15'b000000000000101, 15'b000000000000011, 15'b111111111111111, 15'b000000000000000, 15'b111111111101010, 15'b111111111111111, 15'b000000000000000, 15'b111111111101011, 15'b000000000000000, 15'b000000000000000, 15'b000000000000000, 15'b000000000000000, 15'b111111111010010, 15'b000000000000001, 15'b111111111111111, 15'b111111111111111, 15'b000000000000000, 15'b000000000010000, 15'b111111111111111, 15'b000000000000000, 15'b000000000111010, 15'b000000000101011, 15'b000000000000000, 15'b000000000000000, 15'b111111111100010, 15'b000000000000000, 15'b111111111111111}, 
{15'b000000000001001, 15'b000000000000110, 15'b000000000100000, 15'b111111111100000, 15'b000000000010000, 15'b000000000001111, 15'b000000000000000, 15'b000000000011000, 15'b000000000000001, 15'b111111111111110, 15'b000000000000100, 15'b000000000000000, 15'b111111111111111, 15'b000000000001111, 15'b111111111111111, 15'b111111111111010, 15'b000000000000000, 15'b000000000000100, 15'b111111111111001, 15'b000000000001100, 15'b000000000000100, 15'b111111110110101, 15'b111111111110001, 15'b000000000001011, 15'b111111111111111, 15'b111111110111111, 15'b111111111101111, 15'b111111111111101, 15'b111111111111111, 15'b111111111111000, 15'b000000000000000, 15'b111111111111010}, 
{15'b000000000000000, 15'b111111111111111, 15'b111111111110100, 15'b111111111101010, 15'b000000000000101, 15'b000000000000000, 15'b000000000001100, 15'b111111111111111, 15'b000000000011111, 15'b111111111111111, 15'b000000000000000, 15'b111111111010100, 15'b111111111111111, 15'b000000000010000, 15'b111111111111111, 15'b111111111011110, 15'b000000000000000, 15'b111111111111110, 15'b000000000100001, 15'b111111111111111, 15'b111111111001000, 15'b111111111111111, 15'b000000000100001, 15'b111111111111111, 15'b111111111111111, 15'b000000000010001, 15'b111111111110011, 15'b000000000001000, 15'b000000000000000, 15'b111111111100110, 15'b000000000000000, 15'b000000000000000}, 
{15'b111111111100100, 15'b000000000000000, 15'b000000000000000, 15'b111111111111111, 15'b000000000111111, 15'b111111111110000, 15'b111111111111111, 15'b111111111111111, 15'b111111111111010, 15'b111111111111001, 15'b000000000001000, 15'b000000000010001, 15'b111111111111011, 15'b000000000011111, 15'b000000000000000, 15'b111111111111111, 15'b111111111011011, 15'b111111111111111, 15'b000000000000000, 15'b111111111110101, 15'b000000000000000, 15'b000000000000100, 15'b000000000000001, 15'b111111111111110, 15'b111111111111001, 15'b111111111100110, 15'b111111111011010, 15'b000000000000000, 15'b111111111110001, 15'b000000000000101, 15'b111111111111111, 15'b000000000001001}, 
{15'b111111111001011, 15'b111111111101011, 15'b111111111101100, 15'b000000000000000, 15'b000000001001001, 15'b111111111100011, 15'b000000000000000, 15'b111111111111001, 15'b111111111001011, 15'b000000000010001, 15'b111111111111111, 15'b000000001001000, 15'b000000000000000, 15'b111111111111001, 15'b111111111111111, 15'b000000000000100, 15'b111111111111101, 15'b000000000000000, 15'b111111111111010, 15'b000000000111111, 15'b000000000000100, 15'b111111111111010, 15'b000000000001110, 15'b111111111111111, 15'b111111111111111, 15'b111111111110011, 15'b111111111111010, 15'b111111111000100, 15'b111111111101101, 15'b111111111111111, 15'b111111111111111, 15'b111111111111000}, 
{15'b000000000011100, 15'b111111110011001, 15'b111111110100011, 15'b111111111101010, 15'b000000001010101, 15'b111111111111111, 15'b111111111010011, 15'b000000000100001, 15'b000000000000111, 15'b000000000000000, 15'b000000000011010, 15'b111111111011101, 15'b000000000000000, 15'b000000000000000, 15'b111111111111011, 15'b000000000000010, 15'b111111111110010, 15'b111111110001010, 15'b000000000010101, 15'b000000000101100, 15'b000000000100001, 15'b000000000000000, 15'b000000000000011, 15'b111111111001100, 15'b111111110101111, 15'b111111111111111, 15'b111111111011001, 15'b111111111000101, 15'b111111111100111, 15'b111111110001111, 15'b000000000110101, 15'b000000000110110}, 
{15'b000000000000000, 15'b000000000000000, 15'b000000000000000, 15'b000000000000000, 15'b000000000100001, 15'b111111111101000, 15'b000000000000010, 15'b000000000001001, 15'b111111111010011, 15'b000000000000100, 15'b111111111111111, 15'b111111111111111, 15'b111111111111111, 15'b000000000011110, 15'b000000000000110, 15'b000000000000010, 15'b000000000000111, 15'b000000000101010, 15'b111111111100100, 15'b000000000000000, 15'b111111111101010, 15'b111111111111111, 15'b000000000101000, 15'b000000000000001, 15'b111111111111111, 15'b111111110111000, 15'b111111111111110, 15'b111111111101100, 15'b111111111111000, 15'b000000000000000, 15'b000000000010001, 15'b000000000001101}, 
{15'b111111111111010, 15'b000000000010001, 15'b111111111011001, 15'b000000000000010, 15'b000000000011000, 15'b111111111111010, 15'b111111111111111, 15'b000000000010100, 15'b000000000000000, 15'b111111111111111, 15'b111111111110111, 15'b000000000000000, 15'b000000000000000, 15'b111111111111011, 15'b111111111110000, 15'b111111111110111, 15'b111111111111000, 15'b111111111110111, 15'b111111111110001, 15'b000000000000000, 15'b111111111111111, 15'b111111111111010, 15'b111111111110111, 15'b000000000110010, 15'b000000000000000, 15'b111111111010001, 15'b111111111111110, 15'b000000000001111, 15'b000000000000000, 15'b000000000000000, 15'b000000000100000, 15'b111111111111111}, 
{15'b111111111111111, 15'b000000000000000, 15'b111111111111111, 15'b111111111101100, 15'b111111110010001, 15'b000000000000000, 15'b000000000000000, 15'b111111111111111, 15'b111111110110011, 15'b000000000001010, 15'b111111111110011, 15'b111111111111111, 15'b000000000000000, 15'b111111111010000, 15'b111111111111010, 15'b111111111111111, 15'b000000000000000, 15'b000000000000001, 15'b000000000000100, 15'b000000000101100, 15'b111111111110000, 15'b111111111011001, 15'b000000000000000, 15'b111111111011110, 15'b111111111110011, 15'b111111111100010, 15'b111111111111111, 15'b111111111111110, 15'b111111111111101, 15'b111111111000011, 15'b111111111111011, 15'b000000000011111}, 
{15'b000000000001110, 15'b000000000011100, 15'b111111111111111, 15'b000000000010100, 15'b111111111100101, 15'b111111111110000, 15'b000000000001100, 15'b000000000001000, 15'b111111111111001, 15'b111111111111111, 15'b111111111111111, 15'b111111111111111, 15'b111111111111111, 15'b111111111010110, 15'b111111111111111, 15'b000000000010010, 15'b111111111110001, 15'b000000000000100, 15'b111111111111111, 15'b111111111111111, 15'b000000000011010, 15'b111111111010110, 15'b000000000100011, 15'b000000000000110, 15'b000000000000000, 15'b000000000011011, 15'b000000000000000, 15'b111111111111011, 15'b111111111001111, 15'b111111111110001, 15'b111111111101010, 15'b000000000010110}, 
{15'b000000000000000, 15'b000000000000000, 15'b111111111010001, 15'b111111111111111, 15'b000000000011010, 15'b111111111101101, 15'b111111111111110, 15'b111111111111111, 15'b000000000000010, 15'b000000000000000, 15'b000000000000000, 15'b111111111100101, 15'b000000000001100, 15'b000000000000000, 15'b000000000000000, 15'b000000000000100, 15'b111111111111111, 15'b111111111101100, 15'b000000000000010, 15'b000000000000000, 15'b111111111111011, 15'b111111111111101, 15'b000000000100101, 15'b111111111111111, 15'b000000000000000, 15'b111111111011010, 15'b111111111010110, 15'b000000000011110, 15'b111111111111111, 15'b111111111111111, 15'b000000000000011, 15'b000000000100100}, 
{15'b111111111010100, 15'b111111111111111, 15'b111111111100100, 15'b000000000000000, 15'b111111111010010, 15'b000000000000000, 15'b111111111111111, 15'b111111111110111, 15'b111111110111011, 15'b111111111111100, 15'b000000000000000, 15'b111111111111110, 15'b111111111111111, 15'b000000000000000, 15'b111111111111110, 15'b111111111111001, 15'b111111111101101, 15'b111111111110011, 15'b000000000001000, 15'b111111111111111, 15'b111111111111100, 15'b000000000000000, 15'b000000000101011, 15'b111111111111111, 15'b000000000010011, 15'b000000000001011, 15'b111111111101110, 15'b000000000011011, 15'b111111111111010, 15'b000000000000000, 15'b111111111111111, 15'b000000001001010}, 
{15'b111111111010111, 15'b000000000000011, 15'b000000000000110, 15'b111111111111100, 15'b000000000011111, 15'b111111111011001, 15'b111111111111111, 15'b000000000100001, 15'b000000000010100, 15'b000000000000001, 15'b111111111111111, 15'b111111111110111, 15'b111111111110100, 15'b111111111110111, 15'b111111111111001, 15'b000000000001011, 15'b111111111111111, 15'b000000000000001, 15'b000000000010010, 15'b000000000000000, 15'b000000000000000, 15'b000000000000001, 15'b000000000100000, 15'b000000000000101, 15'b000000000000000, 15'b111111111110010, 15'b111111111111111, 15'b000000000000000, 15'b111111111111110, 15'b111111111111110, 15'b111111111111111, 15'b000000000001000}, 
{15'b111111111111111, 15'b000000000000000, 15'b111111111100100, 15'b111111111110110, 15'b000000000100100, 15'b111111111111111, 15'b111111111110110, 15'b000000000011111, 15'b111111111111001, 15'b000000000100101, 15'b000000000001010, 15'b111111111110000, 15'b000000000000000, 15'b000000000000000, 15'b111111111111110, 15'b000000000000010, 15'b111111111110110, 15'b111111111011110, 15'b000000000100011, 15'b000000000010011, 15'b000000001010001, 15'b000000000011001, 15'b000000000011111, 15'b111111111111111, 15'b000000000000000, 15'b000000000000000, 15'b000000000000111, 15'b000000000001010, 15'b111111111001010, 15'b111111111111111, 15'b111111111111111, 15'b111111111111111}, 
{15'b000000000000000, 15'b111111111110100, 15'b111111111110010, 15'b000000000000000, 15'b111111111100000, 15'b000000000000000, 15'b000000000011000, 15'b000000000001101, 15'b000000000000110, 15'b111111111110011, 15'b000000000000000, 15'b111111111111111, 15'b111111111111111, 15'b111111111111111, 15'b111111111111010, 15'b000000000011001, 15'b111111111111111, 15'b111111111111111, 15'b111111111011001, 15'b000000000000000, 15'b111111111100111, 15'b111111111111111, 15'b000000000000000, 15'b111111111111111, 15'b000000000000001, 15'b000000000000010, 15'b000000000000011, 15'b000000000010001, 15'b111111111110111, 15'b111111111111111, 15'b111111111000110, 15'b000000000001010}, 
{15'b000000000111000, 15'b111111111111110, 15'b000000000001000, 15'b111111111110010, 15'b111111111110101, 15'b000000000000100, 15'b000000000010100, 15'b000000000000000, 15'b000000001000011, 15'b000000000000000, 15'b111111111111101, 15'b000000000000010, 15'b000000000001100, 15'b111111111111111, 15'b000000000000110, 15'b000000000001101, 15'b111111111111111, 15'b111111111000111, 15'b111111111111000, 15'b111111111111111, 15'b000000000001110, 15'b000000000000000, 15'b111111111111111, 15'b000000000001110, 15'b000000000000010, 15'b111111111011110, 15'b111111111110010, 15'b000000000010000, 15'b111111111111100, 15'b000000000100001, 15'b111111111111111, 15'b111111111101001}, 
{15'b000000000000001, 15'b000000000001101, 15'b111111111111111, 15'b111111111111011, 15'b111111111010010, 15'b111111111111111, 15'b000000000000101, 15'b111111111111010, 15'b000000000010101, 15'b111111111111011, 15'b111111111111111, 15'b111111111111011, 15'b111111111111111, 15'b111111111111011, 15'b000000000000000, 15'b000000000101000, 15'b000000000000000, 15'b111111111111111, 15'b111111111111111, 15'b111111111111111, 15'b111111111111111, 15'b111111111111111, 15'b000000000000100, 15'b000000000010000, 15'b000000000000000, 15'b000000000000000, 15'b000000000000100, 15'b111111111111111, 15'b000000000000000, 15'b000000000000010, 15'b000000000000000, 15'b000000000001100}, 
{15'b111111111011000, 15'b000000000010000, 15'b000000000000010, 15'b111111111110010, 15'b111111111001100, 15'b111111111111101, 15'b000000000001000, 15'b111111111001101, 15'b000000001000001, 15'b000000000001001, 15'b000000000000010, 15'b000000000001100, 15'b000000000000101, 15'b000000000000000, 15'b000000000110100, 15'b111111111110101, 15'b000000000000000, 15'b000000000000000, 15'b111111111111111, 15'b000000000000000, 15'b111111111001000, 15'b000000000000010, 15'b000000000010011, 15'b000000000000100, 15'b000000000000100, 15'b111111110101011, 15'b111111111010100, 15'b111111111100001, 15'b000000000000000, 15'b111111111111111, 15'b000000000101001, 15'b111111111100101}, 
{15'b111111111111110, 15'b111111111100111, 15'b111111111110010, 15'b111111111001011, 15'b111111111011110, 15'b000000000101011, 15'b000000000100111, 15'b111111111101010, 15'b000000000000101, 15'b111111111111011, 15'b111111111110011, 15'b111111111011111, 15'b000000000001101, 15'b111111111011011, 15'b000000000011000, 15'b111111111111111, 15'b000000000101010, 15'b111111111111111, 15'b111111111111111, 15'b111111111101110, 15'b111111111111010, 15'b111111111110111, 15'b111111111011101, 15'b000000000001010, 15'b111111111111111, 15'b111111111111111, 15'b111111111100010, 15'b000000000101000, 15'b000000000100011, 15'b111111111110100, 15'b111111110101111, 15'b000000000010010}, 
{15'b000000000000000, 15'b111111111111100, 15'b111111111111111, 15'b111111111110011, 15'b000000000000011, 15'b000000000000001, 15'b000000000001000, 15'b000000000000000, 15'b000000000001111, 15'b111111111111111, 15'b000000000000000, 15'b000000000001100, 15'b000000000000000, 15'b000000000000001, 15'b111111111101111, 15'b111111111110010, 15'b000000000000000, 15'b000000000010111, 15'b000000000000111, 15'b000000000010000, 15'b111111111111101, 15'b111111111101011, 15'b111111111111111, 15'b000000000001001, 15'b111111111111111, 15'b000000000000100, 15'b111111111111111, 15'b000000000001000, 15'b000000000000000, 15'b000000000001010, 15'b111111111001111, 15'b111111111111111}, 
{15'b000000000100111, 15'b111111111111110, 15'b000000000010011, 15'b111111111011000, 15'b111111111100111, 15'b111111111111111, 15'b111111111111111, 15'b000000000000011, 15'b000000000000000, 15'b111111111101111, 15'b000000000000000, 15'b000000000000000, 15'b000000000000000, 15'b000000000000000, 15'b111111111101111, 15'b000000000010010, 15'b111111111111111, 15'b111111111111100, 15'b000000000000000, 15'b000000000001111, 15'b111111111100110, 15'b000000000001110, 15'b000000000010001, 15'b000000000010000, 15'b111111111111111, 15'b000000001000110, 15'b111111111101100, 15'b000000000101110, 15'b111111111111001, 15'b111111111010001, 15'b111111111101001, 15'b000000000010001}, 
{15'b111111110111010, 15'b111111111111100, 15'b111111111101100, 15'b111111111111111, 15'b000000000100001, 15'b111111111101001, 15'b111111111111000, 15'b000000000011110, 15'b000000000001100, 15'b111111111100001, 15'b000000000000000, 15'b111111111111100, 15'b111111111111110, 15'b000000000010001, 15'b111111111100000, 15'b111111111111110, 15'b000000000000000, 15'b111111111111111, 15'b111111111111101, 15'b000000000000000, 15'b111111111100111, 15'b111111111111111, 15'b000000000000000, 15'b111111111010101, 15'b000000000001000, 15'b000000001001111, 15'b000000000101100, 15'b111111111111011, 15'b111111111101011, 15'b111111111000110, 15'b000000000000000, 15'b111111111111001}, 
{15'b000000000000010, 15'b000000000011011, 15'b000000000000010, 15'b111111111101100, 15'b000000000000000, 15'b111111111111100, 15'b000000000000000, 15'b000000000011010, 15'b000000000011011, 15'b111111111101110, 15'b000000000010001, 15'b000000000000011, 15'b111111111111111, 15'b111111111111110, 15'b111111111101011, 15'b000000000100000, 15'b111111111111010, 15'b111111111010110, 15'b000000000001110, 15'b111111111111111, 15'b111111111111111, 15'b000000000001110, 15'b111111111110110, 15'b111111111111111, 15'b111111111111001, 15'b000000000001011, 15'b111111111101110, 15'b000000000010001, 15'b111111111010001, 15'b000000000001010, 15'b111111111111111, 15'b000000000010100}, 
{15'b111111111111010, 15'b000000000000000, 15'b000000000001011, 15'b000000000000000, 15'b111111111111000, 15'b111111111111111, 15'b000000000001101, 15'b111111111111111, 15'b000000000000000, 15'b000000000000000, 15'b000000000000000, 15'b000000000000010, 15'b111111111110010, 15'b000000000000001, 15'b000000000001110, 15'b000000000000101, 15'b000000000001101, 15'b111111111111111, 15'b111111111111111, 15'b000000000010000, 15'b000000000011111, 15'b111111111110011, 15'b000000000000000, 15'b111111111111111, 15'b000000000000001, 15'b111111111000100, 15'b111111111111111, 15'b111111111110110, 15'b111111111111111, 15'b000000001001000, 15'b000000000000000, 15'b111111111100101}, 
{15'b111111111111100, 15'b111111111110000, 15'b111111111111110, 15'b000000000000000, 15'b000000000001011, 15'b111111111111111, 15'b000000000000000, 15'b111111111111101, 15'b000000000001001, 15'b111111111111110, 15'b000000000000000, 15'b000000000000100, 15'b000000000100101, 15'b111111111110010, 15'b000000000000001, 15'b111111110010011, 15'b111111111111110, 15'b111111111111000, 15'b000000000000001, 15'b111111111111001, 15'b000000000001011, 15'b111111111100011, 15'b000000000001110, 15'b000000000001101, 15'b111111111111110, 15'b111111110100100, 15'b111111111100010, 15'b111111111111101, 15'b111111111111101, 15'b000000000110001, 15'b111111111111111, 15'b000000000010011}, 
{15'b000000000000110, 15'b000000000000000, 15'b000000000010110, 15'b111111111110001, 15'b111111111110111, 15'b000000000011110, 15'b111111111101011, 15'b000000000000111, 15'b111111111011000, 15'b000000000000001, 15'b000000000000010, 15'b111111111110101, 15'b000000000000000, 15'b000000000000000, 15'b111111111100111, 15'b000000000110111, 15'b111111111100000, 15'b111111111111110, 15'b000000000001111, 15'b111111111111111, 15'b000000000001000, 15'b111111111000010, 15'b000000000101000, 15'b111111111111111, 15'b111111111110000, 15'b000000000111110, 15'b000000000010010, 15'b111111111101011, 15'b111111111101110, 15'b111111110111011, 15'b111111111111110, 15'b000000000000010}, 
{15'b111111111111111, 15'b000000000000000, 15'b111111111111011, 15'b111111111011101, 15'b111111111111111, 15'b111111111001101, 15'b000000000000000, 15'b000000000100110, 15'b000000000011111, 15'b000000000000010, 15'b000000000000000, 15'b111111111110001, 15'b000000000101010, 15'b111111111111111, 15'b111111111111111, 15'b111111111111111, 15'b000000000110111, 15'b000000000000000, 15'b111111111111010, 15'b111111111111001, 15'b111111111010110, 15'b000000000010000, 15'b000000000000000, 15'b000000000000000, 15'b000000000000100, 15'b111111111110110, 15'b111111111000101, 15'b000000000100011, 15'b111111111000111, 15'b000000000000110, 15'b111111111110101, 15'b000000000000000}, 
{15'b000000000000111, 15'b000000000010111, 15'b000000000000001, 15'b111111111111111, 15'b111111111000101, 15'b000000000000000, 15'b111111111111111, 15'b000000000011111, 15'b000000000100011, 15'b111111111111111, 15'b111111111111111, 15'b111111111111111, 15'b000000000000000, 15'b000000000000000, 15'b000000000000000, 15'b000000000000000, 15'b000000000000000, 15'b111111111111111, 15'b000000000010101, 15'b111111111110010, 15'b111111111001000, 15'b111111111111011, 15'b111111111110011, 15'b111111111110011, 15'b111111111110111, 15'b111111111111111, 15'b111111111110111, 15'b111111111111101, 15'b111111111111110, 15'b000000000010010, 15'b111111111111111, 15'b000000000111011}
};

localparam logic signed [14:0] bias [32] = '{
15'b000000010111100,  // 1.474280834197998
15'b000000001011000,  // 0.6914801001548767
15'b000000010111000,  // 1.4406442642211914
15'b000000010110100,  // 1.408045768737793
15'b000000001111110,  // 0.9864811301231384
15'b000000001101110,  // 0.8636202812194824
15'b111111110110001,  // -0.6153604388237
15'b000000000111101,  // 0.4839226007461548
15'b000000000111110,  // 0.4862793982028961
15'b000000000101111,  // 0.37162142992019653
15'b000000000111010,  // 0.45989668369293213
15'b000000010100110,  // 1.2998151779174805
15'b111111101111101,  // -1.016528844833374
15'b111111111010010,  // -0.35249894857406616
15'b000000000111001,  // 0.44582197070121765
15'b111111111110001,  // -0.1119980737566948
15'b111111111110111,  // -0.06717441976070404
15'b000000000000000,  // 0.00487547367811203
15'b000000000011000,  // 0.1946917623281479
15'b111111110011100,  // -0.7796769738197327
15'b000000001011101,  // 0.7287401556968689
15'b000000011011011,  // 1.714877724647522
15'b111111100110011,  // -1.5971007347106934
15'b000000000001001,  // 0.07393483817577362
15'b000000000101001,  // 0.3225609362125397
15'b000000001101100,  // 0.8453295230865479
15'b000000001110011,  // 0.898597240447998
15'b000000000100000,  // 0.2548799514770508
15'b000000001111100,  // 0.9735668301582336
15'b000000010010000,  // 1.1261906623840332
15'b000000000111001,  // 0.44768181443214417
15'b111111011010000   // -2.3676068782806396
};
endpackage