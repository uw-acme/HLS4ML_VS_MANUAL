// Width: 9
// NFRAC: 4
package dense_4_9_5;

localparam logic signed [8:0] weights [32][5] = '{ 
{9'b111111111, 9'b000000101, 9'b111111011, 9'b000000001, 9'b111111110}, 
{9'b111110111, 9'b111111111, 9'b000000111, 9'b111111111, 9'b000000000}, 
{9'b000000101, 9'b000000011, 9'b111111111, 9'b111111001, 9'b111111100}, 
{9'b111111001, 9'b111111010, 9'b111111110, 9'b000000100, 9'b000000011}, 
{9'b000000001, 9'b000000010, 9'b000000010, 9'b111111111, 9'b111101111}, 
{9'b000000101, 9'b111111001, 9'b000000010, 9'b111111101, 9'b111111101}, 
{9'b111111001, 9'b000000000, 9'b111111111, 9'b000000010, 9'b000000001}, 
{9'b111111111, 9'b000000100, 9'b111111001, 9'b000000010, 9'b000000010}, 
{9'b000000010, 9'b111111101, 9'b000000000, 9'b111111000, 9'b111111100}, 
{9'b111111111, 9'b111111011, 9'b000000010, 9'b000000110, 9'b000000000}, 
{9'b111111101, 9'b111111101, 9'b000000000, 9'b000001001, 9'b111111011}, 
{9'b000000010, 9'b000000011, 9'b111111010, 9'b111111111, 9'b000000001}, 
{9'b000000000, 9'b000000010, 9'b000000000, 9'b111111100, 9'b111110110}, 
{9'b000000010, 9'b000000001, 9'b000000110, 9'b111111110, 9'b111111001}, 
{9'b000000001, 9'b111111111, 9'b111111010, 9'b111111111, 9'b000001000}, 
{9'b111111000, 9'b111111100, 9'b111111100, 9'b000000110, 9'b000000000}, 
{9'b000000101, 9'b111111101, 9'b111111101, 9'b111111100, 9'b111111111}, 
{9'b000000011, 9'b111111111, 9'b111111001, 9'b111111111, 9'b000000001}, 
{9'b000000100, 9'b000000000, 9'b111111100, 9'b000000000, 9'b111111001}, 
{9'b000000011, 9'b111111110, 9'b111111100, 9'b000000011, 9'b000000001}, 
{9'b000000001, 9'b111111111, 9'b000000100, 9'b111111001, 9'b111111111}, 
{9'b000000000, 9'b000000001, 9'b000000111, 9'b111110111, 9'b111110110}, 
{9'b111111110, 9'b000000001, 9'b000000010, 9'b111111010, 9'b000001000}, 
{9'b111111111, 9'b000000010, 9'b000000100, 9'b000000000, 9'b111110110}, 
{9'b111111101, 9'b000000101, 9'b111111100, 9'b000000000, 9'b000000110}, 
{9'b000000000, 9'b000000100, 9'b000000000, 9'b111110100, 9'b000001000}, 
{9'b111111000, 9'b111111100, 9'b000000011, 9'b000000011, 9'b000000011}, 
{9'b000000000, 9'b000000011, 9'b111111111, 9'b111111101, 9'b000000000}, 
{9'b111111110, 9'b000000011, 9'b111110111, 9'b000000010, 9'b111111101}, 
{9'b111111111, 9'b000000010, 9'b111111101, 9'b111111001, 9'b000001001}, 
{9'b000000111, 9'b000000001, 9'b000000101, 9'b111110110, 9'b111111010}, 
{9'b111111111, 9'b111111001, 9'b000000101, 9'b000000001, 9'b000000010}
};

localparam logic signed [8:0] bias [5] = '{
9'b111111111,  // -0.06223141402006149
9'b111111110,  // -0.06270556896924973
9'b111111110,  // -0.07014333456754684
9'b000000001,  // 0.0820775106549263
9'b000000011   // 0.2155742198228836
};
endpackage