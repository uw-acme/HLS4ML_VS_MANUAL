//Width: 37
//Int: 13
package dense_2_gen;

localparam logic signed [36:0] weights [64][32] = '{
{37'b0000000000000010001001101100101010000, 37'b0000000000000000000100001000110101111, 37'b1111111111111110011110110001010010011, 37'b1111111111111111110101001101111110000, 37'b0000000000000010000101101101101000000, 37'b0000000000000000000000000000100110111, 37'b1111111111111110110110000101111101011, 37'b1111111111111111111111111100000000010, 37'b1111111111111101110011110010101100011, 37'b0000000000000000101000110100100011101, 37'b0000000000000000000000000001111100100, 37'b1111111111111111111101000101110110010, 37'b1111111111111111111111110011010111110, 37'b1111111111111110011001100110100010101, 37'b1111111111111111100110000100011001100, 37'b1111111111111101111001111101010001011, 37'b0000000000000000000000000000001111110, 37'b1111111111111111111001010110101101001, 37'b1111111111111110011110011110010111011, 37'b1111111111111110101110111010101001101, 37'b0000000000000000000000000011001001001, 37'b0000000000000000000000000000001111011, 37'b1111111111111111111011111001000100000, 37'b1111111111111111111110100110100010100, 37'b0000000000000000000000000000111010010, 37'b0000000000000000110011011100111101001, 37'b0000000000000011000101101011010100010, 37'b0000000000000001011001101110110111000, 37'b1111111111111111111111110001100100110, 37'b0000000000000000011001111010111111000, 37'b1111111111111100101110011010011001100, 37'b0000000000000000000000001010000100110},
{37'b1111111111111111001100101100101111011, 37'b1111111111111110110000101101010000011, 37'b1111111111111110111001001010111110001, 37'b1111111111111111100011100110100001011, 37'b1111111111111111111101000111101011110, 37'b0000000000000000010110000000111100110, 37'b1111111111111110001101101010111111111, 37'b0000000000000000000010101100010011100, 37'b0000000000000000000010011100000000101, 37'b1111111111111111011111110011111011001, 37'b0000000000000001001111111100000100001, 37'b1111111111111111101001110011100010011, 37'b1111111111111111100001110110110001111, 37'b1111111111111110010000111101110111101, 37'b0000000000000000000011110100100111010, 37'b1111111111111111100111011011110000100, 37'b0000000000000000000110011000100000100, 37'b1111111111111110011100010011101101011, 37'b0000000000000001010111111101100101100, 37'b0000000000000001110101100010110001010, 37'b1111111111111111101111111101111010101, 37'b1111111111111111111101000111010110000, 37'b1111111111111111111111110110111110000, 37'b0000000000000000001100000111011110111, 37'b1111111111111111011011100000010111100, 37'b0000000000000010001100110101100100100, 37'b0000000000000001111110110000010100010, 37'b0000000000000000000100010111110100110, 37'b0000000000000000001110100110110010111, 37'b1111111111111100000110110011001000000, 37'b0000000000000000000011110001000110101, 37'b0000000000000000000000000000001010111},
{37'b0000000000000000100101000110011110010, 37'b1111111111111111000101010001000111010, 37'b1111111111111110111101101001100010001, 37'b1111111111111111101010100110101011111, 37'b1111111111111111011000010111101011100, 37'b1111111111111111010100010101110101001, 37'b1111111111111110100001010101110111110, 37'b0000000000000000000010010010011011111, 37'b1111111111111110111010111000111111000, 37'b0000000000000000000100100100111001100, 37'b0000000000000000000001000100111010010, 37'b1111111111111111010110101100101011101, 37'b0000000000000000101110010010001111011, 37'b1111111111111111011110111110000000100, 37'b1111111111111111111111010011010111111, 37'b1111111111111111101101001101010100110, 37'b0000000000000000000010100001111010100, 37'b0000000000000000110000111001111110101, 37'b0000000000000000011110000000111100100, 37'b0000000000000001110101101011010100100, 37'b0000000000000000010101000010010111101, 37'b1111111111111111010100111100110011101, 37'b0000000000000000000000001100001110000, 37'b0000000000000000010001111001000110101, 37'b1111111111111111110110100110110111110, 37'b0000000000000001101011001010000110100, 37'b0000000000000001001100011000110100111, 37'b0000000000000000110001100110000110111, 37'b1111111111111111111111110010111100011, 37'b1111111111111110110010001000000011100, 37'b1111111111111111111001000100100110001, 37'b0000000000000000110010110110001110000},
{37'b0000000000000001000110101110100000101, 37'b0000000000000000001001110101001100111, 37'b0000000000000000011011000111010011010, 37'b1111111111111111111011000010101000111, 37'b1111111111111011111011010111011001101, 37'b0000000000000000000000000000001011000, 37'b0000000000000000000000001010001111111, 37'b0000000000000001110011110011110011100, 37'b0000000000000001111100001101000001111, 37'b1111111111111111111001001100001110000, 37'b1111111111111111111111111111010000101, 37'b0000000000000000000000000011011000110, 37'b0000000000000000000000001010111110011, 37'b0000000000000000000010100000101000010, 37'b1111111111111111110110101000111010011, 37'b0000000000000001101101111100001011001, 37'b0000000000000000000000000101000001111, 37'b1111111111111111110011011011000111010, 37'b1111111111111111111111111110011010111, 37'b1111111111111110100101110101110001111, 37'b1111111111111111100000101011110001011, 37'b0000000000000000011001010110110100010, 37'b1111111111111111011111100001100010011, 37'b1111111111111111111111110100110101110, 37'b0000000000000000000001111110000100111, 37'b1111111111111111100110000000011000010, 37'b0000000000000000100101011001001110110, 37'b1111111111111111111111111011101110010, 37'b1111111111111111111111111100001101111, 37'b1111111111111111111111111111001010110, 37'b1111111111111110010001110111010110101, 37'b0000000000000010011110110111111010010},
{37'b1111111111111010100010100111001000110, 37'b1111111111111111110011010010110101111, 37'b1111111111111111111101110111111100110, 37'b0000000000000000000010101101111101010, 37'b1111111111111111110010100010111010010, 37'b0000000000000000000011011000100101010, 37'b1111111111111111100110110110000011110, 37'b1111111111111110110011010110110000101, 37'b0000000000000000011011110001101101001, 37'b1111111111111111110101101010111001001, 37'b1111111111111111111001000001111010010, 37'b1111111111111111111111111011100010010, 37'b1111111111111111111111111011010011110, 37'b0000000000000001101011101001010011110, 37'b0000000000000000000000000010111010010, 37'b0000000000000010101000011111101111000, 37'b1111111111111111111111111101011011111, 37'b0000000000000001101111101110100111011, 37'b1111111111111100110011001101011111001, 37'b0000000000000000000000001001110011110, 37'b1111111111111111000110110110111100100, 37'b0000000000000001010110010011110110010, 37'b0000000000000010000100001100111010010, 37'b0000000000000000000000000011101010000, 37'b0000000000000000010111001101111010100, 37'b0000000000000001010011011010101001101, 37'b0000000000000001111010001111101010000, 37'b0000000000000000001000111000000011000, 37'b1111111111111111111101101101100110110, 37'b1111111111111111111111111011001001111, 37'b1111111111111111111000111100001000110, 37'b0000000000000001110011110101101011111},
{37'b0000000000000000011101100010100111001, 37'b1111111111111111111111111010111100101, 37'b0000000000000001001100011010010100000, 37'b1111111111111010110011111111100110100, 37'b1111111111110100111110111001000011110, 37'b1111111111111101001100100101111110111, 37'b0000000000000010110101010111011010000, 37'b1111111111111011000001011111100110101, 37'b1111111111111111111111110101110101111, 37'b1111111111111010100101001100101110010, 37'b1111111111111011111111011110101000011, 37'b1111111111111101010001011000001110100, 37'b0000000000000010110100111010110001000, 37'b1111111111111111111111111110101001101, 37'b1111111111111111111000011001100110001, 37'b0000000000000000000000000001101010000, 37'b1111111111111111111111111111101000111, 37'b1111111111111111111111110010110001111, 37'b1111111111111110111100010011111110101, 37'b1111111111111111111111111100100101011, 37'b1111111111111100000101100001111010101, 37'b0000000000000000000000000000101000010, 37'b0000000000000001011111001101001101101, 37'b1111111111111111111111111101111000100, 37'b0000000000000000001011010001010011000, 37'b0000000000000010001001000100101010110, 37'b0000000000000000011010001111011011000, 37'b1111111111111111111111111111100111111, 37'b1111111111111111111111111100010101111, 37'b0000000000000001101001010000000100011, 37'b1111111111111111101110100001010001100, 37'b0000000000000001100110101100101100110},
{37'b1111111111111111101101100101000000110, 37'b1111111111111110101111011111101001101, 37'b1111111111111110000100010010001111101, 37'b1111111111111111100111111101100010101, 37'b1111111111111101101100010000111010101, 37'b0000000000000000100001110111100001000, 37'b1111111111111110100011110111011111111, 37'b1111111111111110110111010011011111111, 37'b1111111111111100101011101000111000001, 37'b0000000000000000011000110010010001111, 37'b1111111111111111111101011001100111101, 37'b1111111111111110101110100000001000001, 37'b0000000000000000111100111011010010101, 37'b1111111111111111111010110100000101101, 37'b1111111111111111101010110001000000000, 37'b1111111111111011100100100000000110001, 37'b1111111111111111111111111001001111110, 37'b0000000000000000101011000000101110110, 37'b0000000000000001100010001000111101100, 37'b1111111111111110101100111010000111111, 37'b1111111111111110110011001110100001100, 37'b1111111111111111011111111100011011100, 37'b1111111111111111111111010101100010001, 37'b0000000000000000001110001000111110110, 37'b1111111111111111101000101110101101100, 37'b1111111111111010110100001001100011001, 37'b1111111111111101111000010111000100011, 37'b1111111111111111101000111110100010110, 37'b0000000000000000000010111011101010011, 37'b1111111111111111110101000110000000110, 37'b0000000000000000001111101010010001001, 37'b1111111111111111111111101000100000110},
{37'b1111111111111110110001011000000000110, 37'b1111111111111111010001101100111001101, 37'b1111111111111111010111010100011101010, 37'b1111111111111110000110100011001100001, 37'b1111111111111111000100101101011011001, 37'b1111111111111111111111110110010110110, 37'b0000000000000000110101011111001000100, 37'b1111111111111111010111100000111010001, 37'b0000000000000001100110101101110100001, 37'b0000000000000000000000000101000011011, 37'b0000000000000000000000000011111110000, 37'b1111111111111111111111111100000110101, 37'b0000000000000001110000000011111111110, 37'b0000000000000000000000000100100100001, 37'b1111111111111111111111111001110111001, 37'b1111111111111111011011110001011000110, 37'b1111111111111111111111110011111000111, 37'b0000000000000000000000000001111111110, 37'b1111111111111111111111110011001111110, 37'b0000000000000000000000000011100000100, 37'b1111111111111111111111110100101001000, 37'b1111111111111111111111101111001010100, 37'b0000000000000000000000000110100111011, 37'b1111111111111111111111111111010110001, 37'b0000000000000000010110100110000101101, 37'b1111111111111110100011110110111110100, 37'b0000000000000000000111000110000000110, 37'b1111111111111111111111110111110001111, 37'b1111111111111111011011000101111101000, 37'b1111111111111111111111101001101011110, 37'b0000000000000000000000001110110011111, 37'b1111111111111111111111111010111100110},
{37'b1111111111111100001011100011000111110, 37'b1111111111111111100010110000001111100, 37'b1111111111111100111101011000111110000, 37'b0000000000000000111110100111101011000, 37'b0000000000000011111001010100011011100, 37'b1111111111111111111111111111010000101, 37'b1111111111111111110001001000111101100, 37'b0000000000000001111010010100111100100, 37'b1111111111111100011111010110001111101, 37'b1111111111111111101000000101110100001, 37'b0000000000000000000000000011110101111, 37'b1111111111111110011000110110000011110, 37'b1111111111111111111111110100100111010, 37'b0000000000000000100110111111101100100, 37'b1111111111111110011110011101110010001, 37'b0000000000000110000010000000001001001, 37'b1111111111111111111011100111010010010, 37'b0000000000000000010111111100111000010, 37'b0000000000000001101010010111010000001, 37'b0000000000000001111101011000000001011, 37'b0000000000000000000000000110110000001, 37'b1111111111111101010100000100000010001, 37'b0000000000000000000000000111001110101, 37'b0000000000000011010010101110011001111, 37'b1111111111111110100011001111010111000, 37'b0000000000000101100101001100011101001, 37'b1111111111111110110011100101110001101, 37'b1111111111111110010111100111100010100, 37'b1111111111111100001110010111100101011, 37'b1111111111111100010010010110001101001, 37'b0000000000000000000000001001110110000, 37'b0000000000000000011011010110111001000},
{37'b0000000000000000000000000100000111011, 37'b1111111111111111111000000100011111011, 37'b1111111111111111011010001100000001101, 37'b0000000000000000000000000001000011110, 37'b0000000000000010011101111101110110111, 37'b1111111111111111110101101011001011111, 37'b1111111111111111011111011010110101001, 37'b0000000000000000101111000001010010110, 37'b0000000000000000110011111100010001100, 37'b0000000000000000000001110000010011011, 37'b1111111111111111111011101000010110010, 37'b1111111111111111111111110100010100010, 37'b1111111111111111111111111111010010100, 37'b1111111111111111000101110100110000101, 37'b1111111111111111111111111100111000011, 37'b0000000000000000000000001000010010010, 37'b0000000000000000000000000000101000000, 37'b1111111111111111111101011010111110000, 37'b0000000000000000000001000110011100001, 37'b0000000000000000101011011110111101010, 37'b0000000000000000001001110110111000000, 37'b1111111111111111111111111100110000111, 37'b0000000000000000000000000111010000000, 37'b0000000000000000000011101011000001010, 37'b0000000000000000010011101001001111011, 37'b1111111111111110111100011001111111011, 37'b0000000000000000100010110011010100010, 37'b0000000000000001111111010001100110111, 37'b1111111111111111111111111110111010101, 37'b0000000000000000000011001000000100100, 37'b0000000000000000011001011000101111110, 37'b0000000000000000100011100011011011111},
{37'b0000000000000000110001010010100101110, 37'b0000000000000000000000000001100011001, 37'b1111111111111111001011001110001000100, 37'b1111111111111101111111100101000110000, 37'b1111111111111001101001011100100110100, 37'b0000000000000001000100001000000100101, 37'b0000000000000000000000001110100011100, 37'b1111111111111001011000011000100001111, 37'b0000000000000000010010100111101101000, 37'b1111111111111111111111110110101000100, 37'b0000000000000000000001111000100111101, 37'b1111111111111111111111001010101100011, 37'b0000000000000000000101011010001000101, 37'b0000000000000000000000000111110010111, 37'b1111111111111111110110010100101011000, 37'b1111111111111100111100100101110100011, 37'b1111111111111111111111111100001100101, 37'b0000000000000001110000100101001011010, 37'b0000000000000001000000101101010101010, 37'b0000000000000001100001111010110101000, 37'b1111111111111100011110111010010101101, 37'b1111111111111101001001110011001001101, 37'b0000000000000000111101011110101000000, 37'b1111111111111111101110001010100001011, 37'b1111111111111111101000011001011001011, 37'b0000000000000010110111100100001011100, 37'b1111111111111111001110100001010110010, 37'b1111111111111111111111110110110010001, 37'b1111111111111111111111111011101101100, 37'b0000000000000001101100000101111111100, 37'b1111111111111111111111111011001111111, 37'b0000000000000000000011001110000110111},
{37'b1111111111111110011010111110101101000, 37'b1111111111111100000011100101000001101, 37'b0000000000000000000000000000001110001, 37'b1111111111111111111110111010101110111, 37'b0000000000000010101010000001010110000, 37'b1111111111111101110110001011111000011, 37'b1111111111111110001110101001010101101, 37'b0000000000000000111011010110101011110, 37'b1111111111111111111111101100010100110, 37'b0000000000000001001100001010011011110, 37'b0000000000000000100101111001110101000, 37'b1111111111111111011001010000111111011, 37'b0000000000000000000000001000011010100, 37'b0000000000000000000111001111100101001, 37'b1111111111111111110101001001010101100, 37'b1111111111111101111110011100111000111, 37'b0000000000000001011001110100010101010, 37'b0000000000000000001110100110111101000, 37'b0000000000000010011000001100100101010, 37'b0000000000000000101100010011111111101, 37'b0000000000000000000000000001110110101, 37'b1111111111111111101100101001001011101, 37'b0000000000000001000000100010000101100, 37'b1111111111111111010011110000100100110, 37'b1111111111111101100010010010010001001, 37'b1111111111111111111100100100010110010, 37'b0000000000000001011110101110110000100, 37'b1111111111111111111111111001000110100, 37'b0000000000000000000100010100001010100, 37'b1111111111111111001111100001001110110, 37'b0000000000000001000110011001110001010, 37'b0000000000000010001101011100100101110},
{37'b0000000000000000000111110000100001011, 37'b0000000000000000000000000100000011001, 37'b0000000000000001110000010001110010110, 37'b0000000000000000000100010011011010010, 37'b1111111111111111101011001010011100100, 37'b0000000000000001011100011001010101111, 37'b0000000000000000101111001110010011101, 37'b1111111111111111111111110110000000010, 37'b0000000000000000000000011010101010101, 37'b1111111111111110111000001110000101111, 37'b1111111111111111100100000000110000001, 37'b1111111111111110101010010100001101111, 37'b1111111111111111111111111000011110110, 37'b0000000000000000011001110100111110101, 37'b1111111111111111011100101101101100000, 37'b0000000000000110101111101101001010001, 37'b0000000000000000000000001001001111011, 37'b1111111111111111001111110100011001100, 37'b1111111111111110011111011001101010111, 37'b1111111111111111111001001111111001010, 37'b0000000000000001100101101110011001000, 37'b0000000000000001000001100001001000001, 37'b0000000000000000000000000110011000010, 37'b1111111111111111111110101101001011101, 37'b0000000000000001110000011001110111011, 37'b0000000000000010001001010010010000000, 37'b0000000000000011111101100111001110111, 37'b0000000000000000000101010011101000001, 37'b0000000000000000000000000100111011110, 37'b0000000000000000000000001110010010100, 37'b1111111111111111111001111001100101010, 37'b1111111111111111011011011000010011000},
{37'b1111111111111110110000000011100111111, 37'b0000000000000000011000110001011100110, 37'b0000000000000000010100001010100000010, 37'b1111111111111110000001011011010010011, 37'b1111111111111101110110000000001100001, 37'b0000000000000011110000000110010100110, 37'b0000000000000000011001001010101011000, 37'b0000000000000000000000000000011100011, 37'b1111111111111110101101101100011010111, 37'b1111111111111111010010110011001110010, 37'b0000000000000001000010010100001111001, 37'b0000000000000000100100010001010101111, 37'b0000000000000000000000010010101100111, 37'b1111111111111111010111110101110010110, 37'b0000000000000010010010011110001011000, 37'b1111111111111111111111111001000010000, 37'b1111111111111111111001000011000101110, 37'b0000000000000000000000000100111010110, 37'b0000000000000000000110101110000101010, 37'b1111111111111111101000001100101110100, 37'b0000000000000000101000000101111001101, 37'b0000000000000000001000000100101110100, 37'b0000000000000000111010011010011111010, 37'b1111111111111111111111110111111010000, 37'b0000000000000000000001101101111111010, 37'b0000000000000101010000111100100011111, 37'b1111111111111111100011001000100011011, 37'b1111111111111111110100001110100101011, 37'b1111111111111111111111111011100011010, 37'b1111111111111111001000000100101000010, 37'b1111111111111111101011011110111000010, 37'b0000000000000001011010000101111011000},
{37'b0000000000000000011110001011001101101, 37'b0000000000000000100101111110010000001, 37'b0000000000000010100111001010001110010, 37'b1111111111111111101011101001010001100, 37'b0000000000000000110011101100010100100, 37'b0000000000000010110011101001000100110, 37'b0000000000000000000000010110000010111, 37'b1111111111111111110000111100110011001, 37'b0000000000000000111100011010101011000, 37'b1111111111111111000101101101110010111, 37'b1111111111111111111111111100101100010, 37'b1111111111111111000010111111100011110, 37'b0000000000000000000000001010100110000, 37'b0000000000000011001001010100000001000, 37'b1111111111111111110110111101010101111, 37'b0000000000000000000000110100100111101, 37'b0000000000000001111000111010110100000, 37'b0000000000000000000000010101110010000, 37'b0000000000000000000001100000110110101, 37'b1111111111111101011111110101000011001, 37'b1111111111111110000010010010100111001, 37'b1111111111111111101101100001110000011, 37'b1111111111111111111111111111001011110, 37'b1111111111111110110101010011101100011, 37'b1111111111111111101101100001011100001, 37'b1111111111111111010101110010110100101, 37'b1111111111111110011011011100001100100, 37'b1111111111111110010011001110110100100, 37'b0000000000000000001111011000011100001, 37'b0000000000000000111001001001100111110, 37'b1111111111111100110100100111000010000, 37'b0000000000000000000001101010001100110},
{37'b1111111111111101100111001011100011101, 37'b0000000000000000000000000011010101000, 37'b1111111111111111111000011001100000011, 37'b1111111111111111100110100101000100011, 37'b1111111111111111111111111000001001001, 37'b0000000000000001000100010001001110011, 37'b1111111111111111011000011000100111111, 37'b0000000000000010001010110001000111100, 37'b1111111111111101000110000100101000011, 37'b1111111111111111111111101100110100010, 37'b0000000000000000000000000001010100011, 37'b1111111111111111111111111111110010001, 37'b0000000000000000000000001011110001101, 37'b0000000000000000000000000100100101010, 37'b1111111111111111111110000111110001101, 37'b1111111111111111010001100111101101000, 37'b0000000000000000101000100100000010101, 37'b0000000000000001011101110101001000110, 37'b1111111111111111111011001111110010010, 37'b1111111111111101111111010110110111101, 37'b1111111111111111100001111010100111000, 37'b0000000000000000111001010000010100010, 37'b0000000000000000100000010000000100100, 37'b0000000000000000000000001111010111110, 37'b0000000000000000000001100011111001001, 37'b0000000000000000101001110100100101111, 37'b1111111111111110000101011001110001000, 37'b0000000000000000000000000011101111101, 37'b1111111111111111111111111110100111100, 37'b0000000000000000000001101100001111011, 37'b0000000000000000000000010000101100111, 37'b1111111111111110111111100110010110000},
{37'b1111111111111101010011111001101000001, 37'b1111111111111111111101000000110010001, 37'b1111111111111111111110011110101101101, 37'b1111111111111111110111000110100010110, 37'b1111111111111111111101100010000001001, 37'b0000000000000000110110000001000110111, 37'b0000000000000000000011011001000111100, 37'b0000000000000000010001101111110111110, 37'b0000000000000000010011100010010111100, 37'b0000000000000000100000001110010111001, 37'b0000000000000000101000011001000100001, 37'b0000000000000001010010100001100101111, 37'b0000000000000000001101101110000100101, 37'b1111111111111111001110011111000001110, 37'b0000000000000000000000010000001011100, 37'b0000000000000011000011010011111110110, 37'b0000000000000000000000001010011010111, 37'b0000000000000000000000100100101101010, 37'b1111111111111111111110101100111000110, 37'b0000000000000000111000010101110000010, 37'b0000000000000001001000111001001011010, 37'b0000000000000000001111110011010011100, 37'b0000000000000000010101000110010111000, 37'b1111111111111111110000110011001010011, 37'b1111111111111111101111100001110100001, 37'b0000000000000000001101100101010001001, 37'b1111111111111111011101101010010001101, 37'b1111111111111110111111001001110001100, 37'b0000000000000001101011010000101110010, 37'b1111111111111111110000010000011010100, 37'b0000000000000000010000001101010111111, 37'b1111111111111110011111110110011111011},
{37'b0000000000000000000000000100101010001, 37'b1111111111111111111111111110111011110, 37'b0000000000000000010011010010100111000, 37'b0000000000000000000000000100101000001, 37'b0000000000000111010000001111001000111, 37'b1111111111111111111111100111110101110, 37'b0000000000000000000000000000011000111, 37'b1111111111111111111111111111101110011, 37'b0000000000000000111000001001000001000, 37'b1111111111111111011001100010101101110, 37'b0000000000000000000000000000101110010, 37'b0000000000000000000000000010010101010, 37'b0000000000000000000000100100010100010, 37'b0000000000000001000010000111001111010, 37'b0000000000000000000000000001100101100, 37'b1111111111111110110101100100110110000, 37'b1111111111111111111111111101100101110, 37'b1111111111111111011101101100111101111, 37'b0000000000000010100111101001101111100, 37'b0000000000000000000000000111101000111, 37'b1111111111111111111111111111011010011, 37'b1111111111111111111111110110101100100, 37'b0000000000000000000000000011000100000, 37'b1111111111111111111111111111110011010, 37'b0000000000000000000000000001000100111, 37'b0000000000000000100010111111010100011, 37'b0000000000000000000000000001100110111, 37'b0000000000000000000000000001110110001, 37'b1111111111111111111111111111111101000, 37'b1111111111111111111111111011010000011, 37'b0000000000000000000000000111011101111, 37'b0000000000000000010101001101001001111},
{37'b1111111111111111111110010010001111100, 37'b0000000000000000001110110110110010000, 37'b1111111111111111111111100111100100101, 37'b0000000000000000011000100001010100101, 37'b1111111111111111101001010000010101111, 37'b1111111111111111000010111011000001101, 37'b1111111111111111100000000011010011110, 37'b0000000000000010001110001111010100110, 37'b0000000000000000000000001001100101101, 37'b0000000000000000110001100110001111100, 37'b1111111111111111111010010110100010110, 37'b0000000000000000100001001111100100100, 37'b1111111111111111101111000001001010010, 37'b1111111111111110101111010101010100111, 37'b1111111111111110011110011100111001000, 37'b0000000000000000000110101101000001110, 37'b1111111111111111111111111111110000011, 37'b1111111111111111101110001010011011001, 37'b0000000000000000000000000011000000110, 37'b0000000000000000000000001101111111111, 37'b1111111111111111111111101111000011111, 37'b0000000000000000100110110001011010000, 37'b0000000000000000010010010000000000000, 37'b1111111111111110111111100110000001111, 37'b0000000000000000111001001110000000111, 37'b1111111111111110101011110010011100111, 37'b0000000000000000000001000111100011100, 37'b0000000000000000000000000000001110001, 37'b1111111111111110101010001010010000010, 37'b0000000000000000000000000001011010011, 37'b0000000000000000010111010110100001111, 37'b1111111111111111110000000101111110001},
{37'b1111111111111111111010000110110101010, 37'b1111111111111111001101010101100000101, 37'b0000000000000000000000000111011100100, 37'b1111111111111111100001011000110000011, 37'b0000000000000001101110100100011001011, 37'b1111111111111111111111110110101011101, 37'b1111111111111111110101010100101110110, 37'b0000000000000000110110101010001010010, 37'b1111111111111100110111111001110011001, 37'b0000000000000000000000000100001100011, 37'b1111111111111111101100010000100111000, 37'b1111111111111111111110111010010001010, 37'b0000000000000010110011111110000111100, 37'b0000000000000001110101011110000100111, 37'b1111111111111111001101001010110000001, 37'b1111111111111111110101010111100111000, 37'b1111111111111111111111110111101000001, 37'b0000000000000000000000010110001111100, 37'b1111111111111111111111111010011010010, 37'b0000000000000000000000001011001100010, 37'b0000000000000000000000000110001101100, 37'b1111111111111110111010011111010011110, 37'b1111111111111111000011000110100111011, 37'b0000000000000001000011000000010101100, 37'b0000000000000000000000000001011100010, 37'b1111111111111110111001110101001111101, 37'b0000000000000000001100100000110111001, 37'b1111111111111111010110110111010110111, 37'b1111111111111111101110111101111001010, 37'b0000000000000001000101100110001011100, 37'b0000000000000000000000010010011010010, 37'b1111111111111110000001011111101001001},
{37'b0000000000000101000100111110111001001, 37'b0000000000000010101111000101010011110, 37'b1111111111111110000000010110100011011, 37'b0000000000000000000001101010101101010, 37'b1111111111111101001110110100110110101, 37'b0000000000000000000000000010001111011, 37'b0000000000000001110010000101100110000, 37'b0000000000000000001111111011000011100, 37'b0000000000000001110010100101100001111, 37'b1111111111111111111111110110100010111, 37'b1111111111111110110000101111001101011, 37'b1111111111111111010111110011111010101, 37'b0000000000000001001000100100110101100, 37'b0000000000000000001110001010111011101, 37'b1111111111111111001101101110111010100, 37'b0000000000000001000011011100100100010, 37'b0000000000000100010010000010110111100, 37'b1111111111111110111101011011111011010, 37'b1111111111111101101000011001110001100, 37'b0000000000000000000000000010111111001, 37'b1111111111111111110001010100101010000, 37'b1111111111111110100101100100100111001, 37'b1111111111111111111001110011101000010, 37'b1111111111111111111111001110000011110, 37'b0000000000000000101100000000111100110, 37'b1111111111111101000111011110001110101, 37'b0000000000000000101101100001110110010, 37'b1111111111111111111111011100101110001, 37'b0000000000000000000000001010100010010, 37'b0000000000000000110111110101011110000, 37'b1111111111111111110001001111001010010, 37'b0000000000000000011110100000001000000},
{37'b1111111111111111010000100111011110111, 37'b1111111111111110011101101111101011011, 37'b1111111111111111101101011011011011000, 37'b1111111111111110101010010101100100011, 37'b1111111111111111110111001101111101100, 37'b0000000000000000011001001100110110111, 37'b0000000000000000000000000110110011101, 37'b1111111111111111111010001100001001100, 37'b0000000000000000010011010001101010100, 37'b1111111111111111111110001111001101000, 37'b0000000000000000000000000111101110010, 37'b1111111111111110010000111011101011111, 37'b0000000000000000110100001110100101000, 37'b0000000000000000101001001001110010010, 37'b1111111111111111001011100110010111101, 37'b0000000000000011100011000100000011010, 37'b1111111111111111111111111000011101111, 37'b0000000000000000000000000110010011011, 37'b1111111111111111111101111100000100111, 37'b0000000000000000000000000010010100011, 37'b0000000000000010100001110100100000100, 37'b1111111111111100001111000011011100111, 37'b1111111111111111001000100011010001010, 37'b1111111111111111100011010110110000011, 37'b1111111111111111110110011110100101011, 37'b0000000000000001100100111010111111111, 37'b1111111111111111100101001011000110011, 37'b0000000000000000001001000001011000100, 37'b0000000000000011110111111101110000111, 37'b1111111111111011111001100110001100110, 37'b1111111111111101000100000001111001010, 37'b0000000000000000001011011111100010010},
{37'b0000000000000000001000100110111110101, 37'b1111111111111111100001111000010110011, 37'b1111111111111111111111111111101000010, 37'b0000000000000000000000000110111100111, 37'b1111111111111010001111111011000111001, 37'b1111111111111011001001100001110110011, 37'b0000000000000000000000110001011101100, 37'b1111111111111111111111111011010011100, 37'b1111111111111101111000010010101101011, 37'b0000000000000000001100101000000010011, 37'b0000000000000000000000000001010001111, 37'b1111111111111111110001111011001101110, 37'b0000000000000000000000000000101001010, 37'b1111111111111111100010000111111011101, 37'b1111111111111111100101000100001110000, 37'b1111111111111111011100101111111001110, 37'b1111111111111110110100101111011100000, 37'b0000000000000010010000100001011001101, 37'b0000000000000000000000000011100101111, 37'b0000000000000000010111101001100001110, 37'b1111111111111111111111110001111001101, 37'b1111111111111111011011111000100001001, 37'b0000000000000000000000000010011011111, 37'b1111111111111111010011100100011000101, 37'b0000000000000001110000011010000100001, 37'b1111111111111011000001010101001111100, 37'b0000000000000001110000101100101011000, 37'b1111111111111111111111111100001111011, 37'b1111111111111111111101100001010000101, 37'b0000000000000001100110011011101111010, 37'b1111111111111111111111111101000100000, 37'b0000000000000001111000111110101000111},
{37'b1111111111111111111111111010000001011, 37'b0000000000000000000010101001010101111, 37'b1111111111111111101001111010011011111, 37'b0000000000000000100110011110001101010, 37'b0000000000000000011100010101110001010, 37'b1111111111111101010000111011101010101, 37'b0000000000000000000000000111111111100, 37'b0000000000000000100000111110010100001, 37'b0000000000000100101000110000110111100, 37'b1111111111111111111011011010010110010, 37'b0000000000000000000000000000100011001, 37'b0000000000000000011100110110010110001, 37'b0000000000000010110111110010111011001, 37'b1111111111111111101111101111110101010, 37'b0000000000000000000111001010000010000, 37'b0000000000000000110011101110001011011, 37'b1111111111111111111111111100101010001, 37'b0000000000000000001110001110001010111, 37'b1111111111111111111111110110110001100, 37'b0000000000000000000000011110011001011, 37'b1111111111111101110011110111001001010, 37'b0000000000000000010011101000101100101, 37'b0000000000000000100011111110100001000, 37'b0000000000000000001011101000011100010, 37'b1111111111111111111111111011100101001, 37'b0000000000000001101111110000011111001, 37'b0000000000000000000010010011101001001, 37'b0000000000000001000000100010100001101, 37'b1111111111111100101010001100011011111, 37'b0000000000000000110100101000110011001, 37'b0000000000000011001010100101110110010, 37'b0000000000000000000010111001001111111},
{37'b1111111111111101001100010101000110001, 37'b0000000000000001101100000100100011111, 37'b1111111111111101111010101010001001000, 37'b0000000000000000111110111101001111011, 37'b1111111111111111001010000001100101100, 37'b0000000000000000000000001000010111001, 37'b0000000000000011111110110011101011011, 37'b1111111111111110001000110100111000010, 37'b1111111111111101101010111010011000100, 37'b0000000000000001010111101111000011101, 37'b1111111111111110001101111111011110001, 37'b1111111111111111110011111100111001001, 37'b1111111111111111111111100011110101011, 37'b0000000000000010110000001001100011110, 37'b1111111111111111111111001100111101000, 37'b1111111111111101100101100001001000110, 37'b1111111111111111111111111101010001111, 37'b0000000000000011100001101111001000100, 37'b1111111111111100001110110111001110101, 37'b1111111111111111110011100101001100010, 37'b0000000000000010100010000111100100010, 37'b1111111111111101000110010100001000101, 37'b0000000000000000011011001000011101100, 37'b1111111111111111111000010001000101000, 37'b0000000000000010001010111110100011100, 37'b1111111111111011111011100101010001001, 37'b1111111111111101000110010001001001011, 37'b1111111111111110011011100101000000011, 37'b1111111111111111111111111101011011010, 37'b0000000000000000110101000000100100000, 37'b0000000000000000001100110110110110101, 37'b0000000000000001011011010100011111111},
{37'b1111111111111111010001100011001010101, 37'b0000000000000000011010100111110001111, 37'b1111111111111111111111111010110101100, 37'b0000000000000001001100101101000110010, 37'b1111111111111111101100100101101101000, 37'b0000000000000001110100001110100100000, 37'b0000000000000000000001000000111110111, 37'b1111111111111111111010010001101111110, 37'b1111111111111111111110111100100111101, 37'b0000000000000000000000100101011100001, 37'b0000000000000000000000000010011110111, 37'b1111111111111111111111111111100010101, 37'b1111111111111111111111000011111100111, 37'b0000000000000100001010010100111111100, 37'b0000000000000000000110011100110101000, 37'b0000000000000001100000101100000010101, 37'b0000000000000000000000001001001001110, 37'b1111111111111110010011101001100000111, 37'b1111111111111111011000111010110011100, 37'b1111111111111111111111111101010010110, 37'b1111111111111111110111100000110001010, 37'b0000000000000000010101100100010000001, 37'b1111111111111111111111111101101101100, 37'b1111111111111110100001001011110100000, 37'b1111111111111111111111111101100111011, 37'b0000000000000010010111010110010110000, 37'b0000000000000010011110110110000111110, 37'b1111111111111111111111111110010101110, 37'b1111111111111111110111101001111001001, 37'b0000000000000000000000000001001110111, 37'b1111111111111111111111101111100010100, 37'b1111111111111111001110101000001110001},
{37'b1111111111111111010110101001111111011, 37'b0000000000000000000000000010111101010, 37'b0000000000000010001011110000011100011, 37'b0000000000000000000000000010010011100, 37'b0000000000000000000000000011110110100, 37'b1111111111111111000101110111100110000, 37'b0000000000000000000000001011111110100, 37'b1111111111111001000101110000000011101, 37'b0000000000000001101110010110010110101, 37'b0000000000000000000111000010000100000, 37'b0000000000000000001101101011100001111, 37'b1111111111111101000111110000001001100, 37'b0000000000000000000001101111111000111, 37'b1111111111111110111001101001010010000, 37'b1111111111111111101111000000100111010, 37'b0000000000000000000000000101100011111, 37'b0000000000000000001010000011101011000, 37'b0000000000000000000000000110010000100, 37'b0000000000000000111001100011001100110, 37'b0000000000000000000000001001000110110, 37'b1111111111111111111011011101001011100, 37'b0000000000000010101000100100000111100, 37'b0000000000000011000000110001101100100, 37'b1111111111111110001110111001000111011, 37'b1111111111111110110111010001111111001, 37'b0000000000000001111111110001010010100, 37'b1111111111111101100011100001001010010, 37'b0000000000000000001111000001111111000, 37'b1111111111111111111111101100011111111, 37'b1111111111111111111111111100101100001, 37'b1111111111111111111111111001100110111, 37'b0000000000000001011110010010110110101},
{37'b1111111111111111000101111001000001010, 37'b1111111111111111111111101101111000100, 37'b1111111111111110000101100001110111110, 37'b1111111111111110011000100100110100011, 37'b1111111111111111111000111100110010111, 37'b1111111111111110111010111100111110010, 37'b0000000000000000000000000010011101000, 37'b0000000000000000101110101000011100111, 37'b1111111111111110000101010010010101100, 37'b1111111111111111010101010110110000010, 37'b1111111111111111100110100110010010110, 37'b0000000000000000000000001000000001100, 37'b0000000000000000001110010011100001110, 37'b1111111111111111111010111101010111100, 37'b1111111111111111100000110001110101100, 37'b0000000000000000110000111101000111001, 37'b0000000000000001110010000111101001111, 37'b0000000000000001000011001011000000110, 37'b1111111111111110111101000011010011100, 37'b0000000000000000011000111110101101110, 37'b1111111111111111111001111110111100010, 37'b1111111111111111110001011001000000111, 37'b0000000000000000001011100010000001000, 37'b0000000000000000001000001000111111011, 37'b1111111111111111011100011101001000101, 37'b0000000000000000101101100111100010011, 37'b1111111111111111010001100100110000001, 37'b0000000000000000011110101000001011111, 37'b1111111111111111111111111000011000110, 37'b1111111111111101101000110101000111110, 37'b1111111111111111110010100001110111000, 37'b0000000000000001110011001001011001110},
{37'b1111111111111111110010001110011011100, 37'b1111111111111111010101101001000011000, 37'b0000000000000000100111011001100001100, 37'b0000000000000010000001100111000001010, 37'b0000000000000000101011011010000010101, 37'b0000000000000000101010001011111001100, 37'b0000000000000000010111111001110110111, 37'b1111111111111110011000110111111011101, 37'b1111111111111110010110111100000110001, 37'b0000000000000000100011000011111100111, 37'b0000000000000000000110001101101111000, 37'b0000000000000000010110000111010001001, 37'b0000000000000000001011011011110001010, 37'b0000000000000000000010110010000000110, 37'b0000000000000001101001000010111001111, 37'b0000000000000000000011110000010100101, 37'b1111111111111111100100011001010010000, 37'b0000000000000000110100111010101001111, 37'b1111111111111111110000110100110110101, 37'b1111111111111111101101101101010100101, 37'b0000000000000000111000010111011001110, 37'b1111111111111111000000100011101101001, 37'b1111111111111111110010010111001010010, 37'b0000000000000001000001000001100111011, 37'b0000000000000000001011010110110010110, 37'b1111111111111111001001011000010101111, 37'b1111111111111110011010101100110100101, 37'b1111111111111111111001111111001101010, 37'b1111111111111101110001000101001111001, 37'b0000000000000000011110110000010001011, 37'b0000000000000000110100000100011111100, 37'b0000000000000000000000100111010011001},
{37'b1111111111111111111001000010100001000, 37'b1111111111111111110101111001011011010, 37'b1111111111111111111001111011010110000, 37'b1111111111111111101110010000010101011, 37'b1111111111111110111100101001011100011, 37'b1111111111111110111000001011010011011, 37'b0000000000000000100000010101101110100, 37'b0000000000000000000100001111001100100, 37'b1111111111111110100010100101001101000, 37'b0000000000000001010101101100111010010, 37'b1111111111111111110101010110010001101, 37'b1111111111111111111111101100111101001, 37'b1111111111111111000111100110110001110, 37'b0000000000000000000010101011010110100, 37'b0000000000000000001111000111101100010, 37'b1111111111111111100101000100000000110, 37'b1111111111111111110111110111100111100, 37'b1111111111111111101010101001100000011, 37'b1111111111111111010110110111000101000, 37'b0000000000000000000000001001011001100, 37'b1111111111111110111000000111011001111, 37'b0000000000000000110100001011010110001, 37'b1111111111111110010011101110110101011, 37'b0000000000000000000010100011110110010, 37'b0000000000000000010101011111010011011, 37'b0000000000000000111111011101111110100, 37'b0000000000000000001101100111010001100, 37'b0000000000000000000011000100010010100, 37'b0000000000000010010101100000000010100, 37'b0000000000000000011010011011001101100, 37'b0000000000000000000000001000110110110, 37'b0000000000000000101010111011000101100},
{37'b1111111111111111110110000101100100000, 37'b0000000000000010000001011010000010110, 37'b1111111111111111111111111100111010011, 37'b1111111111111111101111001001000010001, 37'b1111111111111110010010100101101111100, 37'b1111111111111111011001100010110100111, 37'b0000000000000011010010101001110110000, 37'b1111111111111010011111001011010101101, 37'b1111111111111101001101000000010110111, 37'b1111111111111110011001110101110110001, 37'b1111111111111110001111101001001011001, 37'b1111111111111101111110001100100110001, 37'b1111111111111111111111101101010100110, 37'b0000000000000011110111111101110001110, 37'b1111111111111111110010100110110110001, 37'b0000000000000000000000000011110100100, 37'b1111111111111110010011111000000000101, 37'b0000000000000011100100001101100100011, 37'b1111111111111100101100101010101011011, 37'b0000000000000000000000000101000100001, 37'b1111111111111111111111110110011011011, 37'b1111111111111101010011110111010010001, 37'b0000000000000000000000000101011000110, 37'b1111111111111111111111111111111111001, 37'b0000000000000000011100110001011001010, 37'b1111111111111111100010100111110101000, 37'b1111111111111110110100010110111010011, 37'b1111111111111111111111111111000110101, 37'b0000000000000001011001011000001001100, 37'b0000000000000000000001101111100000100, 37'b1111111111111111010110111011000110001, 37'b0000000000000000000000011011011110111},
{37'b0000000000000010111100011001111000010, 37'b1111111111111111000110101111101110110, 37'b0000000000000001000011100010111101000, 37'b1111111111111111101111011101101100011, 37'b0000000000000000100111000011111000111, 37'b1111111111111111111110000111010100110, 37'b1111111111111111111110100010000100110, 37'b1111111111111111010000011010110001001, 37'b0000000000000000000000001001100011100, 37'b0000000000000000101111001100011100010, 37'b1111111111111111111111111111011010010, 37'b1111111111111111100001111100011010010, 37'b1111111111111111111111110001011110111, 37'b0000000000000001110101000100001001010, 37'b0000000000000000001001110110111000111, 37'b0000000000000000010100101101001111110, 37'b0000000000000000001100010000010010110, 37'b1111111111111111110011101110000111000, 37'b0000000000000000001010011000100110101, 37'b0000000000000000000000000110000111111, 37'b1111111111111111111011011000101001101, 37'b1111111111111111111111111110100001110, 37'b1111111111111101100011100000101010111, 37'b1111111111111111111111111100111100111, 37'b0000000000000000011101100111010000011, 37'b1111111111111111000100011111001101101, 37'b1111111111111110111010110010110000100, 37'b1111111111111111111111111110000010110, 37'b1111111111111111111111100101100000111, 37'b0000000000000100011101100100111100111, 37'b1111111111111101101101101110011100111, 37'b1111111111111111000100100011000001010},
{37'b1111111111111111101001011100110110001, 37'b1111111111111111001011001000011101000, 37'b1111111111111111011110111111010101010, 37'b0000000000000000010010100101001010110, 37'b0000000000000001000111011011110111110, 37'b1111111111111110111101100001011011111, 37'b1111111111111111111111010101100111011, 37'b1111111111111110001111011100000110000, 37'b0000000000000000011111000110011111011, 37'b0000000000000001000101101001001101100, 37'b1111111111111110010010101111110011111, 37'b1111111111111101111110100100111101100, 37'b0000000000000000001100001101111011010, 37'b1111111111111010100010000111001000011, 37'b1111111111111111011001011011000111010, 37'b1111111111111111000000110001100000011, 37'b1111111111111110011010101111001100010, 37'b1111111111111111111111110100111001000, 37'b0000000000000001000100101111000000100, 37'b0000000000000000000000000001100111100, 37'b1111111111111111101000101000011000101, 37'b1111111111111111101001001010110011111, 37'b0000000000000000000000000001101010000, 37'b0000000000000000000000000011011010000, 37'b1111111111111111100001110011010001010, 37'b1111111111111001111101110010011011101, 37'b1111111111111011100011101011001010110, 37'b1111111111111101110100011110011000110, 37'b0000000000000000011100101000111111010, 37'b0000000000000001101001100111101001010, 37'b1111111111111111111111110111110110110, 37'b0000000000000001111011000010111100011},
{37'b1111111111111111010000110100111100001, 37'b1111111111111110010010000000100011101, 37'b0000000000000001010011110101100111110, 37'b0000000000000000100110001100101101001, 37'b0000000000000000010110001111000111110, 37'b1111111111111111010000111011110000111, 37'b1111111111111111101111010010110101001, 37'b0000000000000000110010011110110101101, 37'b0000000000000100010011111111011100001, 37'b1111111111111110101000010101110001111, 37'b1111111111111111111111111101111110101, 37'b1111111111111111111111111110101001100, 37'b0000000000000000111100001101110100010, 37'b1111111111111111100011111001001100000, 37'b1111111111111111110110110111000001101, 37'b1111111111111111110111011101011101000, 37'b1111111111111111001100110110111101111, 37'b1111111111111111111111100011110100011, 37'b0000000000000000000000000001100001001, 37'b0000000000000001110100000010011000110, 37'b1111111111111110111011111011111110111, 37'b1111111111111111111110011111000101111, 37'b0000000000000001000001110111000010111, 37'b1111111111111111111010110010111001001, 37'b0000000000000000000000000010010100101, 37'b0000000000000100001101011110111011010, 37'b0000000000000010100110000000100111100, 37'b0000000000000000000001101001100100100, 37'b0000000000000000000000001011100001111, 37'b1111111111111100101000100010100110010, 37'b1111111111111111011101000010100001111, 37'b1111111111111111111111111111011000110},
{37'b0000000000000000000111101101011010111, 37'b0000000000000000011000101111110110000, 37'b1111111111111111111000111101011110100, 37'b0000000000000000000000000010011100001, 37'b0000000000000001110110011111101011110, 37'b1111111111111100001000100111101011110, 37'b0000000000000000000000000101001001001, 37'b1111111111111111001111010101110010100, 37'b0000000000000001011111011110001100111, 37'b0000000000000000000000000011001011001, 37'b1111111111111111110110100010001111011, 37'b0000000000000000000000000011010100101, 37'b0000000000000000000000001010110001101, 37'b1111111111111111111111111001110010011, 37'b0000000000000000000010111111000110111, 37'b1111111111111111001000111111001110001, 37'b0000000000000010000100110111011100000, 37'b1111111111111111111101001100011000011, 37'b1111111111111111111000000111000100101, 37'b1111111111111111111111111111111010011, 37'b0000000000000000000000001011000010001, 37'b1111111111111111111100000111110110111, 37'b0000000000000000000000001000011110011, 37'b1111111111111111111111111110010010100, 37'b0000000000000000000110100101011110100, 37'b1111111111111101011101101110010111010, 37'b0000000000000000011010011101010011011, 37'b0000000000000001011101110100001010111, 37'b1111111111111111111110010111010101101, 37'b0000000000000000110000010000000000001, 37'b1111111111111111111111110101100111010, 37'b0000000000000000100110010011011111110},
{37'b1111111111111110011000111111100111111, 37'b0000000000000000000100101011011011000, 37'b1111111111111100001001000001110001101, 37'b0000000000000000000011100010010110000, 37'b1111111111111111100110011011101011000, 37'b1111111111111111101011101000110110000, 37'b1111111111111111111111010111110011011, 37'b1111111111111111010001010111001110011, 37'b1111111111111111101101100110001111101, 37'b1111111111111111011110100011100000111, 37'b0000000000000000011000000101000100111, 37'b0000000000000000001101110001000011000, 37'b1111111111111110100101001110100001101, 37'b0000000000000000000000010001011110011, 37'b1111111111111111111111000011100000111, 37'b1111111111111111111011110110110011101, 37'b0000000000000000100100000101111011110, 37'b1111111111111111110101101000001100011, 37'b1111111111111111110001111001000100111, 37'b1111111111111111110001001001111011101, 37'b1111111111111111111111100110110100100, 37'b0000000000000010001010110000111110110, 37'b1111111111111111111111111110111010010, 37'b0000000000000000000000000010110000001, 37'b1111111111111111111011001101100100000, 37'b0000000000000010100010011101111000101, 37'b0000000000000001100000100111111000000, 37'b0000000000000000010001011010100010101, 37'b1111111111111111001110101001001010101, 37'b1111111111111111111010111011111011110, 37'b0000000000000000100001011001101011010, 37'b0000000000000000011101011110111100001},
{37'b0000000000000000010001011100010000010, 37'b0000000000000000010100000000001110000, 37'b1111111111111111111111111010101010110, 37'b0000000000000000000000001101011001000, 37'b1111111111111100010000000010010000111, 37'b0000000000000000010110010110101100100, 37'b0000000000000000001100101110100101001, 37'b1111111111111111111111110111100001011, 37'b0000000000000000000000010111000010100, 37'b1111111111111110101001001111001011001, 37'b1111111111111111111111111111011010100, 37'b0000000000000000000000000001000011011, 37'b1111111111111110101101101010101001010, 37'b0000000000000000000000000111111011100, 37'b0000000000000000000000001010011011100, 37'b0000000000000000000000001011010000000, 37'b0000000000000000000000000001101101100, 37'b1111111111111101001001110101110000010, 37'b0000000000000000000100111000101111011, 37'b1111111111111111111111101111001110100, 37'b1111111111111111111111110011001001001, 37'b0000000000000000000000000101010000010, 37'b0000000000000001000010000001110011100, 37'b1111111111111111111111111100110001111, 37'b0000000000000000000000000100100110010, 37'b0000000000000011101001011010010011000, 37'b0000000000000010101110001010011101110, 37'b0000000000000000000000000101111001010, 37'b0000000000000000000000000101100010011, 37'b1111111111111110001000011010111110001, 37'b0000000000000000000000001100011001010, 37'b1111111111111111111111111101100001100},
{37'b0000000000000000100110110011000100110, 37'b0000000000000000011011000000010011110, 37'b0000000000000010000001100110000010100, 37'b1111111111111110000000111000010011100, 37'b0000000000000001000011110000101110000, 37'b0000000000000000111100110010101111101, 37'b0000000000000000000011001101001001111, 37'b0000000000000001100010001101111110001, 37'b0000000000000000000110000110000111000, 37'b1111111111111111111001110111101101001, 37'b0000000000000000010011000111000111100, 37'b0000000000000000000010111101110111111, 37'b1111111111111111111111101110101110111, 37'b0000000000000000111101110000011101000, 37'b1111111111111111111101001000001111000, 37'b1111111111111111101011101111101100101, 37'b0000000000000000000000010111101111110, 37'b0000000000000000010000010010010110101, 37'b1111111111111111100111010100100000101, 37'b0000000000000000110010100011101011101, 37'b0000000000000000010000101000111111110, 37'b1111111111111011010110110100001010100, 37'b1111111111111111000101011010011110101, 37'b0000000000000000101110110001110000010, 37'b1111111111111111111111111111011110111, 37'b1111111111111011111101011110001100100, 37'b1111111111111110111111011011101100010, 37'b1111111111111111110100001101101101001, 37'b1111111111111111111111101010000111101, 37'b1111111111111111100010110000010111010, 37'b0000000000000000000000000001101011101, 37'b1111111111111111101011101111111111110},
{37'b0000000000000000000000111100000010110, 37'b1111111111111111111111111100010010011, 37'b1111111111111111010001001010101010010, 37'b1111111111111110101001110110000100001, 37'b0000000000000000010101011111011100010, 37'b0000000000000000000000000110111011101, 37'b0000000000000000110000110011101001011, 37'b1111111111111111111101000100011010111, 37'b0000000000000001111111110010100011001, 37'b1111111111111111111101111100001011001, 37'b0000000000000000000000000011110001011, 37'b1111111111111101010000001010001110111, 37'b1111111111111111111111110011011011110, 37'b0000000000000001000000011110111111111, 37'b1111111111111111111111111001100000111, 37'b1111111111111101111010100011110011111, 37'b0000000000000000000000000001111011001, 37'b1111111111111111111010001101001110101, 37'b0000000000000010000110100111100000110, 37'b1111111111111111111111111110101111110, 37'b1111111111111100100000011111000000110, 37'b1111111111111111111111111100001111011, 37'b0000000000000010000100000111000001101, 37'b1111111111111111111111111101011111111, 37'b1111111111111111111111111101000001000, 37'b0000000000000001000111000111011000001, 37'b1111111111111111001111111101100010001, 37'b0000000000000000100011011010101001000, 37'b0000000000000000000000000111111101110, 37'b1111111111111110011000110110111011000, 37'b0000000000000000000000000011011000111, 37'b0000000000000000000001010000011000011},
{37'b1111111111111110010001010011111110010, 37'b0000000000000000000000100101110110010, 37'b0000000000000000000000010001010001100, 37'b1111111111111111111100111011101100001, 37'b0000000000000011111101110100110100010, 37'b1111111111111111000000011010111101001, 37'b1111111111111111111101001001011100101, 37'b1111111111111111111100010000000111000, 37'b1111111111111111101001000110101001011, 37'b1111111111111111100110001100110000110, 37'b0000000000000000100001011000001011010, 37'b0000000000000001000100000001100000110, 37'b1111111111111111101101001010100010101, 37'b0000000000000001111111110000010001100, 37'b0000000000000000000000000101011011111, 37'b1111111111111111111111110011111101101, 37'b1111111111111101101110100011011110101, 37'b1111111111111111111111101101101001101, 37'b0000000000000000000000001110111001101, 37'b1111111111111111010111001111010100111, 37'b0000000000000000000001000100100011101, 37'b0000000000000000010011000110110111010, 37'b0000000000000000000110110110101110100, 37'b1111111111111111111011010100101100100, 37'b1111111111111111100101111111111110001, 37'b1111111111111110011000001000010000011, 37'b1111111111111101101000100010011000001, 37'b0000000000000000000000001000000010011, 37'b1111111111111111000110000000110010110, 37'b0000000000000000010100011000000101100, 37'b1111111111111111111111110101110100111, 37'b0000000000000000100110101110001100000},
{37'b1111111111111100101100011101101011111, 37'b1111111111111110101111111011001001101, 37'b1111111111111110110000000010101110011, 37'b0000000000000000000000000010111111000, 37'b0000000000000100100100011110111101101, 37'b1111111111111110001110000011110000101, 37'b0000000000000000000000000010001000011, 37'b1111111111111111100100010000110110111, 37'b1111111111111100101110001010110101111, 37'b0000000000000001000110111011101111100, 37'b1111111111111111111111111111010100100, 37'b0000000000000100100010011000010100101, 37'b0000000000000000000000001110101110110, 37'b1111111111111111100111101110001001111, 37'b1111111111111111111111110111111101000, 37'b0000000000000000010000001110100000111, 37'b1111111111111111110110011110110111100, 37'b0000000000000000000000001110001100011, 37'b1111111111111111101000001011110001010, 37'b0000000000000011111101101001010010010, 37'b0000000000000000010011110110101111011, 37'b1111111111111111101010101001101101100, 37'b0000000000000000111000000101000110110, 37'b1111111111111111111111110110100110000, 37'b1111111111111111111111111110101110110, 37'b1111111111111111001110001111101101101, 37'b1111111111111111101000000001010001101, 37'b1111111111111100010000011100111110011, 37'b1111111111111110110110000100000000101, 37'b1111111111111111111111111110011001110, 37'b1111111111111111111111011110000111000, 37'b1111111111111111100001111110010010100},
{37'b0000000000000001110011101010001110001, 37'b1111111111111001100110101001011100011, 37'b1111111111111010001101000110110001100, 37'b1111111111111110101000111000110110101, 37'b0000000000000101010110101101010111001, 37'b1111111111111111111111111110100001101, 37'b1111111111111101001110100000110000111, 37'b0000000000000010000111100110111010000, 37'b0000000000000000011110011000011010101, 37'b0000000000000000000000011101001011100, 37'b0000000000000001101010101110101110101, 37'b1111111111111101110101000010000111001, 37'b0000000000000000000000011100101111100, 37'b0000000000000000000010001100100010111, 37'b1111111111111111101111111111101111010, 37'b0000000000000000001001001110110000111, 37'b1111111111111111001010110111100110111, 37'b1111111111111000101000001101011000101, 37'b0000000000000001010101111011010110011, 37'b0000000000000010110000100100000001000, 37'b0000000000000010000111101111111111000, 37'b0000000000000000000001010110100110011, 37'b0000000000000000001110111000001100000, 37'b1111111111111100110001101110100011010, 37'b1111111111111010111100000011001010010, 37'b1111111111111111111101011110011100011, 37'b1111111111111101100110100000001110111, 37'b1111111111111100010101100101010110100, 37'b1111111111111110011100001101011010110, 37'b1111111111111000111110111101110110000, 37'b0000000000000011010110101000000110110, 37'b0000000000000011011011110010000001000},
{37'b0000000000000000000000001000001100110, 37'b0000000000000000000000010100010001110, 37'b0000000000000000000001001001101011101, 37'b0000000000000000000000000110101001101, 37'b0000000000000010000100100100111110100, 37'b1111111111111110100000010000111101011, 37'b0000000000000000001001000111111110010, 37'b0000000000000000100101010110111100000, 37'b1111111111111101001101010100100110010, 37'b0000000000000000010010110011011011100, 37'b1111111111111111111101101100011010011, 37'b1111111111111111111111100000110100110, 37'b1111111111111111111111111010000001000, 37'b0000000000000001111010101011010100110, 37'b0000000000000000011010100100101101000, 37'b0000000000000000001011001000001001101, 37'b0000000000000000011111101001011101100, 37'b0000000000000010101010101000010100000, 37'b1111111111111110010000001001111111000, 37'b0000000000000000000000000011111010100, 37'b1111111111111110101011111001010100111, 37'b1111111111111111111111110110101100000, 37'b0000000000000010100001000111100101110, 37'b0000000000000000000100001010110001000, 37'b1111111111111111111110100011111001110, 37'b1111111111111011100000101110000001001, 37'b1111111111111111111011010011111111101, 37'b1111111111111110110000111110011010011, 37'b1111111111111111100000110011001011000, 37'b0000000000000000000001110100010011100, 37'b0000000000000001000101001010001001010, 37'b0000000000000000110101000101110101110},
{37'b1111111111111111101001110110011110111, 37'b0000000000000001000100100100101101100, 37'b1111111111111101100100011100100011110, 37'b0000000000000000001010100101110011011, 37'b0000000000000001100011001001100011110, 37'b1111111111111111101011110000000010101, 37'b1111111111111111111101101000010110001, 37'b0000000000000001010011100111100110001, 37'b0000000000000000000000001000110100010, 37'b1111111111111111111111111001101000000, 37'b1111111111111111011110100001001111011, 37'b0000000000000000000000000000111010100, 37'b0000000000000000000000001100100110110, 37'b1111111111111111101110011111000110010, 37'b1111111111111111000001101100011111010, 37'b1111111111111111011110000011001000101, 37'b1111111111111111100011001001000001101, 37'b1111111111111111011111110100110111011, 37'b1111111111111111000111110010010111100, 37'b0000000000000000000000000011111011101, 37'b1111111111111111111111110110101001010, 37'b1111111111111111101001000111010000011, 37'b1111111111111111011101111000101111010, 37'b0000000000000011001011101011001100010, 37'b0000000000000000000000000000111011111, 37'b1111111111111101000111101100010001000, 37'b1111111111111111111011101011001101101, 37'b0000000000000000111111000101010101101, 37'b0000000000000000000000001110000101100, 37'b0000000000000000000000000000000111110, 37'b0000000000000010000000011111110110001, 37'b1111111111111111111111110010011010010},
{37'b1111111111111111111111111100101011101, 37'b0000000000000000000010000110100010111, 37'b1111111111111111111111110100101101101, 37'b1111111111111110110000000000010110101, 37'b1111111111111001000111100001101111101, 37'b0000000000000000000000011110001011001, 37'b0000000000000000000000001010010111011, 37'b1111111111111111111100101011001111110, 37'b1111111111111011001101000010010011100, 37'b0000000000000000101001110001100010010, 37'b1111111111111111001101110011000111110, 37'b1111111111111111111111111110000101110, 37'b0000000000000000000000001111100010011, 37'b1111111111111101000010100101111111011, 37'b1111111111111111101000100011111111111, 37'b1111111111111111111111110111001011001, 37'b0000000000000000000000101100100010110, 37'b0000000000000000000100001111001011100, 37'b0000000000000000010010100101010011100, 37'b0000000000000010110000110001011111000, 37'b1111111111111111000010110000001111011, 37'b1111111111111101100110111001111101100, 37'b0000000000000000000000000011101111110, 37'b1111111111111101111011111110100000011, 37'b1111111111111111001101011111000000010, 37'b1111111111111110001001100011010110111, 37'b1111111111111111111100001101111111011, 37'b1111111111111111111001100110000001111, 37'b1111111111111111110110101101000001011, 37'b1111111111111100001110110010011101011, 37'b1111111111111111101110100011101011111, 37'b0000000000000001111100000010101010011},
{37'b0000000000000000111001111110101100100, 37'b0000000000000001110000001110101100110, 37'b1111111111111111111110111111000010011, 37'b0000000000000001010001100100011010011, 37'b1111111111111110010100000000010000110, 37'b1111111111111111000000010001110000001, 37'b0000000000000000110000111101101000001, 37'b0000000000000000100011001010010001001, 37'b1111111111111111100111111010000100111, 37'b1111111111111111111111111100000111100, 37'b1111111111111111111111111100000110111, 37'b1111111111111111111111111001001001101, 37'b1111111111111111111111110110000011110, 37'b1111111111111101011011111110110010101, 37'b1111111111111111111111111101100111110, 37'b0000000000000001001001110110001010000, 37'b1111111111111111000101011101111101001, 37'b0000000000000000010001110101100011011, 37'b1111111111111111111111010100101100000, 37'b1111111111111111111111011110011110100, 37'b0000000000000001101010001100000111110, 37'b1111111111111101011000100001110110101, 37'b0000000000000010001111110010100100000, 37'b0000000000000000011000010100111110001, 37'b0000000000000000000000001000100111011, 37'b0000000000000001101100011111011000100, 37'b0000000000000000000001100111111110010, 37'b1111111111111111101101100001000001101, 37'b1111111111111100111101001011111010111, 37'b1111111111111111000111111111000011101, 37'b1111111111111110101000110101010011110, 37'b0000000000000001011010111010010011010},
{37'b0000000000000000000000000000110100001, 37'b0000000000000000000011101100001000001, 37'b1111111111111101000100101011010111111, 37'b1111111111111111111110110001000010010, 37'b0000000000000001101001110101111110011, 37'b1111111111111110110111100001001010001, 37'b1111111111111111111001110100110001001, 37'b1111111111111111111111111101101000010, 37'b0000000000000000001010011011010111111, 37'b0000000000000000000000000001100000010, 37'b0000000000000000000000000000110100110, 37'b1111111111111110010111101010000100000, 37'b0000000000000000110001001010001100011, 37'b0000000000000000000011000110100111010, 37'b0000000000000000000000000101001001100, 37'b0000000000000000010011001010110000101, 37'b1111111111111111111111110101011100101, 37'b1111111111111110110011110111001100011, 37'b0000000000000000001001001010011101110, 37'b0000000000000000000000000101101110010, 37'b1111111111111111101110011011010010100, 37'b1111111111111111110100110001110100000, 37'b0000000000000010010111101101101000111, 37'b1111111111111111111111111101000101010, 37'b0000000000000000000000000010000100000, 37'b1111111111111101101010001010001110011, 37'b1111111111111101011000101001110011111, 37'b0000000000000001111011100111010010010, 37'b1111111111111111111111010110110101101, 37'b1111111111111111111111110100100111011, 37'b0000000000000000001110001011101110010, 37'b0000000000000010010000101101110110011},
{37'b1111111111111101010001100010000011100, 37'b1111111111111111111111111110001011111, 37'b1111111111111110010011000110010000001, 37'b0000000000000000000010001100000010110, 37'b1111111111111101001011000101011010000, 37'b0000000000000000000000000000000111001, 37'b1111111111111111111111110111101111001, 37'b1111111111111111011110100010000001010, 37'b1111111111111011101111011101111100000, 37'b1111111111111111110010110100111010001, 37'b0000000000000000000000000011001101010, 37'b1111111111111111111011110000011110100, 37'b1111111111111111111111110101000101101, 37'b0000000000000000000000000010110011110, 37'b1111111111111111111011100111011001101, 37'b1111111111111111100110100010011011111, 37'b1111111111111110110100011111001101001, 37'b1111111111111111001111001010111010111, 37'b0000000000000000100001111001111100100, 37'b1111111111111111111110110001110010001, 37'b1111111111111111110011000011011000100, 37'b0000000000000000000000000010011101011, 37'b0000000000000010101100011000000000111, 37'b1111111111111111111111111011100001110, 37'b0000000000000001001100100000111010001, 37'b0000000000000000101110111100110111110, 37'b1111111111111110111001100011001101111, 37'b0000000000000001101101001100111100010, 37'b1111111111111111101000100100110000110, 37'b0000000000000000000000000001011110111, 37'b1111111111111111111111011010110001110, 37'b0000000000000100101010000000100111111},
{37'b1111111111111101011111001111011010001, 37'b0000000000000000001111001101110011101, 37'b0000000000000000011001111100001110100, 37'b1111111111111111110001101000001111001, 37'b0000000000000001111101000010110010000, 37'b1111111111111101100101010000001100111, 37'b1111111111111111111100011011000001101, 37'b0000000000000010000111111111100000001, 37'b0000000000000001010001100100000100010, 37'b0000000000000000000100101101110111101, 37'b1111111111111111111111111100010100110, 37'b1111111111111111011100111101110100101, 37'b1111111111111111010010001100010111111, 37'b1111111111111111011110111000010010001, 37'b1111111111111111100110100101101110100, 37'b0000000000000000101110001100011101100, 37'b1111111111111111111111111100000111111, 37'b0000000000000000000100001001010000100, 37'b0000000000000001001000010111011000110, 37'b0000000000000000000000000010111000001, 37'b0000000000000000000000000011110011011, 37'b0000000000000000000111101001111000010, 37'b0000000000000010000001000001111111010, 37'b0000000000000000010111011010001101001, 37'b0000000000000000000011011011001100001, 37'b1111111111111111001000111010010001101, 37'b1111111111111111111111111100110101101, 37'b0000000000000000000000000000110110101, 37'b1111111111111111111000110000000111010, 37'b1111111111111111111001110100011100001, 37'b1111111111111111111111110110000100111, 37'b0000000000000000100010100110100010010},
{37'b1111111111111111111111111010100111010, 37'b0000000000000000000001111110101111001, 37'b1111111111111110010011011101101101000, 37'b1111111111111111011001110110101110111, 37'b0000000000000010010000011101111100010, 37'b1111111111111111111111110100111001001, 37'b1111111111111111011000010111111110111, 37'b0000000000000001111101001011011010101, 37'b1111111111111111100100111000111111011, 37'b0000000000000010010101010100110101100, 37'b0000000000000000101011110010110011110, 37'b1111111111111111000010011101110010001, 37'b0000000000000000000000010010011000111, 37'b0000000000000000000001110011100110100, 37'b1111111111111111111000011111010101111, 37'b0000000000000000001010111000100110000, 37'b1111111111111111011000100011000010110, 37'b1111111111111101111001001100011001000, 37'b0000000000000010001110010011111100000, 37'b0000000000000001001111100010001110100, 37'b0000000000000101000100111110000101110, 37'b0000000000000001100110110000010010011, 37'b0000000000000001111111000001010010000, 37'b1111111111111111111111111000101000000, 37'b0000000000000000000000000001001110011, 37'b0000000000000000000000000001101001101, 37'b0000000000000000011101010111100001111, 37'b0000000000000000101000100100110100100, 37'b1111111111111100101000111111110001000, 37'b1111111111111111111111111001011010110, 37'b1111111111111111111101011000100011101, 37'b1111111111111111111100101001001101111},
{37'b0000000000000000000000010001001000011, 37'b1111111111111111010011001001001000100, 37'b1111111111111111001010111111010010001, 37'b0000000000000000000000000001111110100, 37'b1111111111111110000011010000000000100, 37'b0000000000000000000000000010100111010, 37'b0000000000000001100010000001100010011, 37'b0000000000000000110111111001000111011, 37'b0000000000000000011011001100011100111, 37'b1111111111111111001101011101000110011, 37'b0000000000000000000000000010011110011, 37'b1111111111111111111111111110010001111, 37'b1111111111111111111111111000100011010, 37'b1111111111111111111111111010101001010, 37'b1111111111111111101010001010100111011, 37'b0000000000000001100111011100011000011, 37'b1111111111111111111111111110101101110, 37'b1111111111111111111111101111010010101, 37'b1111111111111101100101001101100101001, 37'b0000000000000000000000000101111000110, 37'b1111111111111110011101011111101110000, 37'b1111111111111111111111011111011110101, 37'b0000000000000000000000000101111101011, 37'b1111111111111111111101111001100100100, 37'b0000000000000000000111101110000000011, 37'b0000000000000000001000111011110100011, 37'b0000000000000000001110010011010110000, 37'b0000000000000001000110110111001100010, 37'b1111111111111111011110101110000010010, 37'b1111111111111111111100000101101010001, 37'b1111111111111100011010010011000111011, 37'b0000000000000000101000010111001111010},
{37'b0000000000000011100010001101011000110, 37'b1111111111111111111011100011100000000, 37'b0000000000000000100001111010000010111, 37'b1111111111111111001010011001010011001, 37'b1111111111111111010100010010011011100, 37'b0000000000000000010001000101101000101, 37'b0000000000000001010010000010010001110, 37'b0000000000000000000000000010110011101, 37'b0000000000000100001101110101100101101, 37'b0000000000000000000000001010101010101, 37'b1111111111111111110101000010010111101, 37'b0000000000000000001001101011001000010, 37'b0000000000000000110000001010100101001, 37'b1111111111111111111110101011000010100, 37'b0000000000000000011011010000010000000, 37'b0000000000000000110100111001110001111, 37'b1111111111111111111101110011111010010, 37'b1111111111111100011100000101010000111, 37'b1111111111111111100011001000000010101, 37'b1111111111111111111111001001111000111, 37'b0000000000000000111011100010101010110, 37'b0000000000000000000000110111111010000, 37'b1111111111111111111111110000010000001, 37'b0000000000000000111001100110000000011, 37'b0000000000000000001001001100101011001, 37'b1111111111111101111001000010010010101, 37'b1111111111111111001011011010111001001, 37'b0000000000000001000011101100111001110, 37'b1111111111111111110001100010011000101, 37'b0000000000000010000100001001100111001, 37'b1111111111111111111111011100010001001, 37'b1111111111111110100100011111010101110},
{37'b0000000000000000000110101001000001010, 37'b0000000000000000110100001011010001011, 37'b1111111111111111111111111110100100111, 37'b1111111111111111101100001011101101011, 37'b1111111111111101001011010010001100011, 37'b1111111111111111111111110010110101011, 37'b0000000000000000010111100100001011110, 37'b1111111111111111101000011011110011110, 37'b0000000000000001010100011011110010010, 37'b1111111111111111101110100000100100111, 37'b1111111111111111111111100100111001100, 37'b1111111111111111101110111001101010011, 37'b1111111111111111111111111000000001111, 37'b1111111111111111101101000011100001000, 37'b0000000000000000000000000010111100110, 37'b0000000000000010100000010010110110000, 37'b0000000000000000000000000010001111001, 37'b1111111111111111111111000111110000011, 37'b1111111111111111111111111000010010001, 37'b1111111111111111111111111010101001000, 37'b1111111111111111111111111000010000001, 37'b1111111111111111111111110010101001000, 37'b0000000000000000010001011101110010011, 37'b0000000000000001000000011101110111110, 37'b0000000000000000000000000000100011111, 37'b0000000000000000000010001000011010000, 37'b0000000000000000010000100101010000010, 37'b1111111111111111111111101110010111100, 37'b0000000000000000000000000010110111000, 37'b0000000000000000001010011100100100110, 37'b0000000000000000000000110001010100101, 37'b0000000000000000110001100100001101100},
{37'b1111111111111101100001111000000100001, 37'b0000000000000001000010101100111011110, 37'b0000000000000000001001001101001110101, 37'b1111111111111111001010001111101100000, 37'b1111111111111100110011100100100011001, 37'b1111111111111111110110101000000000010, 37'b0000000000000000100010010011000010110, 37'b1111111111111100110100100000110000100, 37'b0000000000000100000101111010111101001, 37'b0000000000000000100100101100000011111, 37'b0000000000000000001000000000100011011, 37'b0000000000000000110000010000110011100, 37'b0000000000000000010110101101011100100, 37'b0000000000000000000000010110101110101, 37'b0000000000000011010000110011011010010, 37'b1111111111111111010100111011011111100, 37'b0000000000000000000010101010100101111, 37'b0000000000000000000000000011010010010, 37'b1111111111111111111100100100011011110, 37'b0000000000000000000001111011101111100, 37'b1111111111111100100010111100001011111, 37'b0000000000000000001000101011010010111, 37'b0000000000000001001110010010011100010, 37'b0000000000000000010011001111100100001, 37'b0000000000000000010010011110110011110, 37'b1111111111111010101111111110101000100, 37'b1111111111111101010001011110111101001, 37'b1111111111111110000100110010000111101, 37'b0000000000000000000001010111101011101, 37'b1111111111111111111111000110001110001, 37'b0000000000000010100110110111111010011, 37'b1111111111111110010111001011000101001},
{37'b1111111111111111111001011011001001110, 37'b1111111111111110011100011111111101010, 37'b1111111111111111001011000100011001101, 37'b1111111111111100101110110001010010111, 37'b1111111111111101111010110010101111011, 37'b0000000000000010101100001001000011111, 37'b0000000000000010011110101010010100110, 37'b1111111111111110101000111010011111010, 37'b0000000000000000010101010011001100000, 37'b1111111111111111101100001001110111010, 37'b1111111111111111001111111010010111011, 37'b1111111111111101111111010011010001100, 37'b0000000000000000110100110011011000111, 37'b1111111111111101101110100000100011101, 37'b0000000000000001100000101000011100110, 37'b1111111111111111111111110101000100110, 37'b0000000000000010101011111110000101000, 37'b1111111111111111111111111111111011101, 37'b1111111111111111111100000000001110110, 37'b1111111111111110111010101100101001101, 37'b1111111111111111101010101101100111010, 37'b1111111111111111011110111111011111011, 37'b1111111111111101110111111111110000101, 37'b0000000000000000101010001011100111001, 37'b1111111111111111111111111100100010110, 37'b1111111111111111111100110000110101001, 37'b1111111111111110001011001011010000001, 37'b0000000000000010100001001101110010011, 37'b0000000000000010001110111000111110110, 37'b1111111111111111010001101100001010110, 37'b1111111111111010111101001011011010111, 37'b0000000000000001001001001000110101110},
{37'b0000000000000000000000001100100101011, 37'b1111111111111111110010111010101110111, 37'b1111111111111111111111111001000100100, 37'b1111111111111111001110001111001000011, 37'b0000000000000000001110100101011100000, 37'b0000000000000000000100101010110000100, 37'b0000000000000000100011101011010000101, 37'b0000000000000000000010111100111010111, 37'b0000000000000000111100010111000111011, 37'b1111111111111111111111100001011001110, 37'b0000000000000000000000000000000100101, 37'b0000000000000000110000110110110110100, 37'b0000000000000000000000111100011001100, 37'b0000000000000000000110010000101000100, 37'b1111111111111110111100001111111111011, 37'b1111111111111111001000110110111100010, 37'b0000000000000000000000000010100011000, 37'b0000000000000001011101000011110011000, 37'b0000000000000000011101000101110000101, 37'b0000000000000001000000011000100111000, 37'b1111111111111111110111100010010110101, 37'b1111111111111110101110001010011001101, 37'b1111111111111111111111111010001011110, 37'b0000000000000000100110000010101100010, 37'b1111111111111111111111111011100000000, 37'b0000000000000000010000100100111111100, 37'b1111111111111111111101100010001010001, 37'b0000000000000000100010100100110010100, 37'b0000000000000000000000000110111111001, 37'b0000000000000000101010100101010010111, 37'b1111111111111100111101101101011001111, 37'b1111111111111111111111111101101100100},
{37'b0000000000000010011110111011110110010, 37'b1111111111111111111011011000110011001, 37'b0000000000000001001100110000111010110, 37'b1111111111111101100011101110001101011, 37'b1111111111111110011101001000111101011, 37'b1111111111111111111111111101001010110, 37'b1111111111111111111111111011101011000, 37'b0000000000000000001110000000010111101, 37'b0000000000000000000001001100000010111, 37'b1111111111111110111111100001101001110, 37'b0000000000000000000000000000101011110, 37'b0000000000000000000001000000011101011, 37'b0000000000000000000000000001000000100, 37'b0000000000000000000000001010111101111, 37'b1111111111111110111101111001011001011, 37'b0000000000000001001001000001100111110, 37'b1111111111111111111111001011011111000, 37'b1111111111111111110000001011110000001, 37'b0000000000000000000000000100110001101, 37'b0000000000000000111101011101100001100, 37'b1111111111111110011001001100100001001, 37'b0000000000000000111011011111100100010, 37'b0000000000000001000111101111000100011, 37'b0000000000000001000010000010001001110, 37'b1111111111111111111111111110100111101, 37'b0000000000000100011010010111000000001, 37'b1111111111111110110001100110110110110, 37'b0000000000000010111010000100011111011, 37'b1111111111111111100101100111111100000, 37'b1111111111111101000111010110011010111, 37'b1111111111111110100111001111000011010, 37'b0000000000000001000111011000010100000},
{37'b1111111111111011101001111011101000001, 37'b1111111111111111110010010101000110111, 37'b1111111111111110110001001001010001011, 37'b1111111111111111111111111110100011001, 37'b0000000000000010000101100001010000100, 37'b1111111111111110100100100110010010001, 37'b1111111111111111100001010101001001100, 37'b0000000000000001111001111110111101001, 37'b0000000000000000110000011011101100010, 37'b1111111111111110000110001010000010111, 37'b0000000000000000000000000100110000110, 37'b1111111111111111110001100110001101010, 37'b1111111111111111111010111110111100000, 37'b0000000000000001000110011010110100101, 37'b1111111111111110000010001101110110101, 37'b1111111111111111111010010001010110100, 37'b0000000000000000000000000001111001100, 37'b1111111111111111111111101010110101000, 37'b1111111111111111110111110010011011000, 37'b0000000000000000000000000011110011101, 37'b1111111111111110011110101011001110111, 37'b1111111111111111111111111001101111100, 37'b0000000000000000000000000010100111111, 37'b1111111111111101010111111001011011011, 37'b0000000000000000100011111100011011010, 37'b0000000000000100111101010111100100100, 37'b0000000000000010110001000100100010000, 37'b1111111111111111101101101010101001001, 37'b1111111111111110101101110010011001000, 37'b1111111111111100011010010010111000011, 37'b0000000000000000000000001010111101100, 37'b1111111111111111100111000000111111010},
{37'b0000000000000000001010111110000110011, 37'b0000000000000001101101011011101010110, 37'b0000000000000000001010111001000111000, 37'b1111111111111110110010101000010011101, 37'b0000000000000000000010010110110101001, 37'b1111111111111111110010111110111110101, 37'b0000000000000000000000000110010010111, 37'b0000000000000001101010101110111010010, 37'b0000000000000001101110000011001101101, 37'b1111111111111110111011100101000001110, 37'b0000000000000001000111111011111010001, 37'b0000000000000000001100010011010001111, 37'b1111111111111111111111111101100011100, 37'b1111111111111111111000101101100000001, 37'b1111111111111110101110101101001000000, 37'b0000000000000010000001100000100001100, 37'b1111111111111111101010010010111000100, 37'b1111111111111101011010100100101000011, 37'b0000000000000000111010100011000001111, 37'b1111111111111111111111111010111110111, 37'b1111111111111111111111111001001100010, 37'b0000000000000000111011110101010010001, 37'b1111111111111111011001111100101110011, 37'b1111111111111111111101100010001010100, 37'b1111111111111111100101100101011111101, 37'b0000000000000000101101001000010001110, 37'b1111111111111110111000001011001010001, 37'b0000000000000001000100101011110000000, 37'b1111111111111101000101110000101111111, 37'b0000000000000000101001001100111110011, 37'b1111111111111111111111110001101011101, 37'b0000000000000001010000001101100101100},
{37'b1111111111111111101010000010101111101, 37'b0000000000000000000000010011010001000, 37'b0000000000000000101101100101011000000, 37'b0000000000000000000000000011011101101, 37'b1111111111111111100000110000011100111, 37'b1111111111111111111110100010100111111, 37'b0000000000000000110100100011010011001, 37'b1111111111111111111111111110100111101, 37'b0000000000000000000000000111111100100, 37'b0000000000000000000010100110100100001, 37'b0000000000000000000000000101010000110, 37'b0000000000000000001010001101000001111, 37'b1111111111111111001001100101011110110, 37'b0000000000000000000101010101010111000, 37'b0000000000000000111000101101010000110, 37'b0000000000000000010111111011001101010, 37'b0000000000000000110110000010111011110, 37'b1111111111111111111111101110111101110, 37'b1111111111111111111111010100011000011, 37'b0000000000000001000001100010000000010, 37'b0000000000000001111110101010110110001, 37'b1111111111111111001101111011001001101, 37'b0000000000000000000000000010000010110, 37'b1111111111111111111110111101001011111, 37'b0000000000000000000101110110101001111, 37'b1111111111111100010011111110101110011, 37'b1111111111111111111111100101010111001, 37'b1111111111111111011011110001000110000, 37'b1111111111111111111111111000110101011, 37'b0000000000000100100001000100001001101, 37'b0000000000000000000000001000110101011, 37'b1111111111111110010110100100111001101},
{37'b1111111111111111110010010000011000101, 37'b1111111111111111000010111001101100001, 37'b1111111111111111111011011111011001101, 37'b0000000000000000000011100101110001100, 37'b0000000000000000101110011100110001011, 37'b1111111111111111111111111100100000100, 37'b0000000000000000000000000111110101000, 37'b1111111111111111110100001001110100110, 37'b0000000000000000100100001011110100010, 37'b1111111111111111111011110011010000100, 37'b0000000000000000000000000100111011000, 37'b0000000000000000010000001101110111111, 37'b0000000000000010010111000011101111010, 37'b1111111111111111001011110010100110001, 37'b0000000000000000000110011101001011100, 37'b1111111111111001001101101101011110000, 37'b1111111111111111111010010010110111010, 37'b1111111111111111100001000010001110010, 37'b0000000000000000000100000110000001111, 37'b1111111111111111100110011100100111010, 37'b0000000000000000101111000111000011111, 37'b1111111111111110001101010000001111100, 37'b0000000000000000111010011101001011011, 37'b0000000000000000110101111110101110101, 37'b1111111111111111111001010010011100000, 37'b1111111111111010010011111101000011101, 37'b1111111111111110001010111111101001001, 37'b1111111111111111110100110100101010000, 37'b1111111111111111110110100111001110100, 37'b0000000000000011000111111101101101010, 37'b1111111111111111111101000001110000101, 37'b0000000000000001001110111001110110010},
{37'b0000000000000000011000000011100010010, 37'b0000000000000000000000000101010010010, 37'b0000000000000001011001001011100001110, 37'b1111111111111111000101111011111100010, 37'b1111111111111111011100110011100001101, 37'b0000000000000001111001110010111101011, 37'b1111111111111110101110001000110100011, 37'b0000000000000000011101011100001000011, 37'b1111111111111101100001100101010101011, 37'b0000000000000000000100011111010111000, 37'b0000000000000000001000100101011011010, 37'b1111111111111111010101000011110011101, 37'b0000000000000000000000010001101001111, 37'b0000000000000000000000000000000001000, 37'b1111111111111110011111110100001100100, 37'b0000000000000011011101011011111101111, 37'b1111111111111110000001101010111000010, 37'b1111111111111111111001111001111000001, 37'b0000000000000000111100110110011001010, 37'b1111111111111111111111111011010110111, 37'b0000000000000000100011011111001001101, 37'b1111111111111100001010101100100100001, 37'b0000000000000010100000010110001101000, 37'b1111111111111111111111111110000110100, 37'b1111111111111111000000100110010001010, 37'b0000000000000011111000001001101101110, 37'b0000000000000001001010110010001001010, 37'b1111111111111110101111001110001101001, 37'b1111111111111110111011001011110111010, 37'b1111111111111011101100111110111111110, 37'b1111111111111111111010110010010010100, 37'b0000000000000000001000001000101101100},
{37'b1111111111111111111111111111000001110, 37'b0000000000000000000011010111100111011, 37'b1111111111111111101110001101100110010, 37'b1111111111111101110110110011101111111, 37'b1111111111111111111111110101101001011, 37'b1111111111111100110111000101101000001, 37'b0000000000000000000000001001010011011, 37'b0000000000000010011011011100101110010, 37'b0000000000000001111101000100110011110, 37'b0000000000000000001001101010110011011, 37'b0000000000000000000000000000101111100, 37'b1111111111111111000111100111001110101, 37'b0000000000000010101010000010110100100, 37'b1111111111111111111111111110110010100, 37'b1111111111111111111111110101110110101, 37'b1111111111111111111111110010011101110, 37'b0000000000000011011110001011001001001, 37'b0000000000000000000000110100001000010, 37'b1111111111111111101011101010001000101, 37'b1111111111111111100101110111101001101, 37'b1111111111111101011011001101101100011, 37'b0000000000000001000011011000000001000, 37'b0000000000000000000000000000010101110, 37'b0000000000000000000000000001101101000, 37'b0000000000000000010000001100010110101, 37'b1111111111111111011011100101100111110, 37'b1111111111111100010100001011010011111, 37'b0000000000000010001101010000110111100, 37'b1111111111111100011100111111001101010, 37'b0000000000000000011010001011100011000, 37'b1111111111111111010111100101111011111, 37'b0000000000000000000000000000010000101},
{37'b0000000000000000011111011000011111100, 37'b0000000000000001011111011101010000011, 37'b0000000000000000000100111100001010000, 37'b1111111111111111111110011110100000010, 37'b1111111111111100010100110111111001000, 37'b0000000000000000000000011101110011100, 37'b1111111111111111111111111110100100101, 37'b0000000000000001111100000011011111011, 37'b0000000000000010001101110110000100100, 37'b1111111111111111111111111010010000101, 37'b1111111111111111111111111011010111010, 37'b1111111111111111111111010111111111101, 37'b0000000000000000000000000101011110001, 37'b0000000000000000000001000011101010110, 37'b0000000000000000000000000000000000000, 37'b0000000000000000000000000110110111011, 37'b0000000000000000000000001110100001011, 37'b1111111111111111111111101011011111111, 37'b0000000000000001010111000000011110101, 37'b1111111111111111001011010010011110110, 37'b1111111111111100100010110101001100010, 37'b1111111111111111101111000010000100100, 37'b1111111111111111001101011000000101111, 37'b1111111111111111001111111101111011011, 37'b1111111111111111011100100011011100111, 37'b1111111111111111111111100010000100101, 37'b1111111111111111011111110011000010010, 37'b1111111111111111110100110010101110111, 37'b1111111111111111111010101011011000000, 37'b0000000000000001001000011010110000111, 37'b1111111111111111111111110101101111100, 37'b0000000000000011101101010010101110111}
};
localparam logic signed [36:0] bias [32] = '{
37'b0000000000001011110010110101001111000,
37'b0000000000000101100010000010011010111,
37'b0000000000001011100001100111000010000,
37'b0000000000001011010000111010110110000,
37'b0000000000000111111001000101000000111,
37'b0000000000000110111010001011000111000,
37'b1111111111111011000100111011110111101,
37'b0000000000000011110111110001001011010,
37'b0000000000000011111000111110011001110,
37'b0000000000000010111110010001010010101,
37'b0000000000000011101011011101111001010,
37'b0000000000001010011001100000010110000,
37'b1111111111110111110111100010011000100,
37'b1111111111111101001011100001010100001,
37'b0000000000000011100100010000101100100,
37'b1111111111111111000110101010000011000,
37'b1111111111111111011101100110110101000,
37'b0000000000000000000010011111110000101,
37'b0000000000000001100011101011101010010,
37'b1111111111111001110000110011100010111,
37'b0000000000000101110101000111010110111,
37'b0000000000001101101110000001000111010,
37'b1111111111110011001110010010001101000,
37'b0000000000000000100101110110101100101,
37'b0000000000000010100101001001101011010,
37'b0000000000000110110000110011110000100,
37'b0000000000000111001100000101001111000,
37'b0000000000000010000010011111111010000,
37'b0000000000000111110010011101110101101,
37'b0000000000001001000000100111000001000,
37'b0000000000000011100101001101101000110,
37'b1111111111101101000011110010010000100
};
endpackage