// Width: 16
// NFRAC: 6
package dense_2_16_6;

localparam logic signed [15:0] weights [64][32] = '{ 
{16'b0000000000010001, 16'b0000000000000000, 16'b1111111111110011, 16'b1111111111111110, 16'b0000000000010000, 16'b0000000000000000, 16'b1111111111110110, 16'b1111111111111111, 16'b1111111111101110, 16'b0000000000000101, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111110011, 16'b1111111111111100, 16'b1111111111101111, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111110011, 16'b1111111111110101, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000110, 16'b0000000000011000, 16'b0000000000001011, 16'b1111111111111111, 16'b0000000000000011, 16'b1111111111100101, 16'b0000000000000000}, 
{16'b1111111111111001, 16'b1111111111110110, 16'b1111111111110111, 16'b1111111111111100, 16'b1111111111111111, 16'b0000000000000010, 16'b1111111111110001, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111011, 16'b0000000000001001, 16'b1111111111111101, 16'b1111111111111100, 16'b1111111111110010, 16'b0000000000000000, 16'b1111111111111100, 16'b0000000000000000, 16'b1111111111110011, 16'b0000000000001010, 16'b0000000000001110, 16'b1111111111111101, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000001, 16'b1111111111111011, 16'b0000000000010001, 16'b0000000000001111, 16'b0000000000000000, 16'b0000000000000001, 16'b1111111111100000, 16'b0000000000000000, 16'b0000000000000000}, 
{16'b0000000000000100, 16'b1111111111111000, 16'b1111111111110111, 16'b1111111111111101, 16'b1111111111111011, 16'b1111111111111010, 16'b1111111111110100, 16'b0000000000000000, 16'b1111111111110111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111010, 16'b0000000000000101, 16'b1111111111111011, 16'b1111111111111111, 16'b1111111111111101, 16'b0000000000000000, 16'b0000000000000110, 16'b0000000000000011, 16'b0000000000001110, 16'b0000000000000010, 16'b1111111111111010, 16'b0000000000000000, 16'b0000000000000010, 16'b1111111111111110, 16'b0000000000001101, 16'b0000000000001001, 16'b0000000000000110, 16'b1111111111111111, 16'b1111111111110110, 16'b1111111111111111, 16'b0000000000000110}, 
{16'b0000000000001000, 16'b0000000000000001, 16'b0000000000000011, 16'b1111111111111111, 16'b1111111111011111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000001110, 16'b0000000000001111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111110, 16'b0000000000001101, 16'b0000000000000000, 16'b1111111111111110, 16'b1111111111111111, 16'b1111111111110100, 16'b1111111111111100, 16'b0000000000000011, 16'b1111111111111011, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111100, 16'b0000000000000100, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111110010, 16'b0000000000010011}, 
{16'b1111111111010100, 16'b1111111111111110, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111110, 16'b0000000000000000, 16'b1111111111111100, 16'b1111111111110110, 16'b0000000000000011, 16'b1111111111111110, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000001101, 16'b0000000000000000, 16'b0000000000010101, 16'b1111111111111111, 16'b0000000000001101, 16'b1111111111100110, 16'b0000000000000000, 16'b1111111111111000, 16'b0000000000001010, 16'b0000000000010000, 16'b0000000000000000, 16'b0000000000000010, 16'b0000000000001010, 16'b0000000000001111, 16'b0000000000000001, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000001110}, 
{16'b0000000000000011, 16'b1111111111111111, 16'b0000000000001001, 16'b1111111111010110, 16'b1111111110100111, 16'b1111111111101001, 16'b0000000000010110, 16'b1111111111011000, 16'b1111111111111111, 16'b1111111111010100, 16'b1111111111011111, 16'b1111111111101010, 16'b0000000000010110, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111110111, 16'b1111111111111111, 16'b1111111111100000, 16'b0000000000000000, 16'b0000000000001011, 16'b1111111111111111, 16'b0000000000000001, 16'b0000000000010001, 16'b0000000000000011, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000001101, 16'b1111111111111101, 16'b0000000000001100}, 
{16'b1111111111111101, 16'b1111111111110101, 16'b1111111111110000, 16'b1111111111111100, 16'b1111111111101101, 16'b0000000000000100, 16'b1111111111110100, 16'b1111111111110110, 16'b1111111111100101, 16'b0000000000000011, 16'b1111111111111111, 16'b1111111111110101, 16'b0000000000000111, 16'b1111111111111111, 16'b1111111111111101, 16'b1111111111011100, 16'b1111111111111111, 16'b0000000000000101, 16'b0000000000001100, 16'b1111111111110101, 16'b1111111111110110, 16'b1111111111111011, 16'b1111111111111111, 16'b0000000000000001, 16'b1111111111111101, 16'b1111111111010110, 16'b1111111111101111, 16'b1111111111111101, 16'b0000000000000000, 16'b1111111111111110, 16'b0000000000000001, 16'b1111111111111111}, 
{16'b1111111111110110, 16'b1111111111111010, 16'b1111111111111010, 16'b1111111111110000, 16'b1111111111111000, 16'b1111111111111111, 16'b0000000000000110, 16'b1111111111111010, 16'b0000000000001100, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000001110, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111011, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000010, 16'b1111111111110100, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111011, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111}, 
{16'b1111111111100001, 16'b1111111111111100, 16'b1111111111100111, 16'b0000000000000111, 16'b0000000000011111, 16'b1111111111111111, 16'b1111111111111110, 16'b0000000000001111, 16'b1111111111100011, 16'b1111111111111101, 16'b0000000000000000, 16'b1111111111110011, 16'b1111111111111111, 16'b0000000000000100, 16'b1111111111110011, 16'b0000000000110000, 16'b1111111111111111, 16'b0000000000000010, 16'b0000000000001101, 16'b0000000000001111, 16'b0000000000000000, 16'b1111111111101010, 16'b0000000000000000, 16'b0000000000011010, 16'b1111111111110100, 16'b0000000000101100, 16'b1111111111110110, 16'b1111111111110010, 16'b1111111111100001, 16'b1111111111100010, 16'b0000000000000000, 16'b0000000000000011}, 
{16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111011, 16'b0000000000000000, 16'b0000000000010011, 16'b1111111111111110, 16'b1111111111111011, 16'b0000000000000101, 16'b0000000000000110, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000101, 16'b0000000000000001, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000010, 16'b1111111111110111, 16'b0000000000000100, 16'b0000000000001111, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000011, 16'b0000000000000100}, 
{16'b0000000000000110, 16'b0000000000000000, 16'b1111111111111001, 16'b1111111111101111, 16'b1111111111001101, 16'b0000000000001000, 16'b0000000000000000, 16'b1111111111001011, 16'b0000000000000010, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111110, 16'b1111111111100111, 16'b1111111111111111, 16'b0000000000001110, 16'b0000000000001000, 16'b0000000000001100, 16'b1111111111100011, 16'b1111111111101001, 16'b0000000000000111, 16'b1111111111111101, 16'b1111111111111101, 16'b0000000000010110, 16'b1111111111111001, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000001101, 16'b1111111111111111, 16'b0000000000000000}, 
{16'b1111111111110011, 16'b1111111111100000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000010101, 16'b1111111111101110, 16'b1111111111110001, 16'b0000000000000111, 16'b1111111111111111, 16'b0000000000001001, 16'b0000000000000100, 16'b1111111111111011, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111110, 16'b1111111111101111, 16'b0000000000001011, 16'b0000000000000001, 16'b0000000000010011, 16'b0000000000000101, 16'b0000000000000000, 16'b1111111111111101, 16'b0000000000001000, 16'b1111111111111010, 16'b1111111111101100, 16'b1111111111111111, 16'b0000000000001011, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111001, 16'b0000000000001000, 16'b0000000000010001}, 
{16'b0000000000000000, 16'b0000000000000000, 16'b0000000000001110, 16'b0000000000000000, 16'b1111111111111101, 16'b0000000000001011, 16'b0000000000000101, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111110111, 16'b1111111111111100, 16'b1111111111110101, 16'b1111111111111111, 16'b0000000000000011, 16'b1111111111111011, 16'b0000000000110101, 16'b0000000000000000, 16'b1111111111111001, 16'b1111111111110011, 16'b1111111111111111, 16'b0000000000001100, 16'b0000000000001000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000001110, 16'b0000000000010001, 16'b0000000000011111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111011}, 
{16'b1111111111110110, 16'b0000000000000011, 16'b0000000000000010, 16'b1111111111110000, 16'b1111111111101110, 16'b0000000000011110, 16'b0000000000000011, 16'b0000000000000000, 16'b1111111111110101, 16'b1111111111111010, 16'b0000000000001000, 16'b0000000000000100, 16'b0000000000000000, 16'b1111111111111010, 16'b0000000000010010, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111101, 16'b0000000000000101, 16'b0000000000000001, 16'b0000000000000111, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000101010, 16'b1111111111111100, 16'b1111111111111110, 16'b1111111111111111, 16'b1111111111111001, 16'b1111111111111101, 16'b0000000000001011}, 
{16'b0000000000000011, 16'b0000000000000100, 16'b0000000000010100, 16'b1111111111111101, 16'b0000000000000110, 16'b0000000000010110, 16'b0000000000000000, 16'b1111111111111110, 16'b0000000000000111, 16'b1111111111111000, 16'b1111111111111111, 16'b1111111111111000, 16'b0000000000000000, 16'b0000000000011001, 16'b1111111111111110, 16'b0000000000000000, 16'b0000000000001111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111101011, 16'b1111111111110000, 16'b1111111111111101, 16'b1111111111111111, 16'b1111111111110110, 16'b1111111111111101, 16'b1111111111111010, 16'b1111111111110011, 16'b1111111111110010, 16'b0000000000000001, 16'b0000000000000111, 16'b1111111111100110, 16'b0000000000000000}, 
{16'b1111111111101100, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111100, 16'b1111111111111111, 16'b0000000000001000, 16'b1111111111111011, 16'b0000000000010001, 16'b1111111111101000, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111010, 16'b0000000000000101, 16'b0000000000001011, 16'b1111111111111111, 16'b1111111111101111, 16'b1111111111111100, 16'b0000000000000111, 16'b0000000000000100, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000101, 16'b1111111111110000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111110111}, 
{16'b1111111111101010, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111110, 16'b1111111111111111, 16'b0000000000000110, 16'b0000000000000000, 16'b0000000000000010, 16'b0000000000000010, 16'b0000000000000100, 16'b0000000000000101, 16'b0000000000001010, 16'b0000000000000001, 16'b1111111111111001, 16'b0000000000000000, 16'b0000000000011000, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000111, 16'b0000000000001001, 16'b0000000000000001, 16'b0000000000000010, 16'b1111111111111110, 16'b1111111111111101, 16'b0000000000000001, 16'b1111111111111011, 16'b1111111111110111, 16'b0000000000001101, 16'b1111111111111110, 16'b0000000000000010, 16'b1111111111110011}, 
{16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000010, 16'b0000000000000000, 16'b0000000000111010, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000111, 16'b1111111111111011, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000001000, 16'b0000000000000000, 16'b1111111111110110, 16'b1111111111111111, 16'b1111111111111011, 16'b0000000000010100, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000100, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000010}, 
{16'b1111111111111111, 16'b0000000000000001, 16'b1111111111111111, 16'b0000000000000011, 16'b1111111111111101, 16'b1111111111111000, 16'b1111111111111100, 16'b0000000000010001, 16'b0000000000000000, 16'b0000000000000110, 16'b1111111111111111, 16'b0000000000000100, 16'b1111111111111101, 16'b1111111111110101, 16'b1111111111110011, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111101, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000100, 16'b0000000000000010, 16'b1111111111110111, 16'b0000000000000111, 16'b1111111111110101, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111110101, 16'b0000000000000000, 16'b0000000000000010, 16'b1111111111111110}, 
{16'b1111111111111111, 16'b1111111111111001, 16'b0000000000000000, 16'b1111111111111100, 16'b0000000000001101, 16'b1111111111111111, 16'b1111111111111110, 16'b0000000000000110, 16'b1111111111100110, 16'b0000000000000000, 16'b1111111111111101, 16'b1111111111111111, 16'b0000000000010110, 16'b0000000000001110, 16'b1111111111111001, 16'b1111111111111110, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111110111, 16'b1111111111111000, 16'b0000000000001000, 16'b0000000000000000, 16'b1111111111110111, 16'b0000000000000001, 16'b1111111111111010, 16'b1111111111111101, 16'b0000000000001000, 16'b0000000000000000, 16'b1111111111110000}, 
{16'b0000000000101000, 16'b0000000000010101, 16'b1111111111110000, 16'b0000000000000000, 16'b1111111111101001, 16'b0000000000000000, 16'b0000000000001110, 16'b0000000000000001, 16'b0000000000001110, 16'b1111111111111111, 16'b1111111111110110, 16'b1111111111111010, 16'b0000000000001001, 16'b0000000000000001, 16'b1111111111111001, 16'b0000000000001000, 16'b0000000000100010, 16'b1111111111110111, 16'b1111111111101101, 16'b0000000000000000, 16'b1111111111111110, 16'b1111111111110100, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000101, 16'b1111111111101000, 16'b0000000000000101, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000110, 16'b1111111111111110, 16'b0000000000000011}, 
{16'b1111111111111010, 16'b1111111111110011, 16'b1111111111111101, 16'b1111111111110101, 16'b1111111111111110, 16'b0000000000000011, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000010, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111110010, 16'b0000000000000110, 16'b0000000000000101, 16'b1111111111111001, 16'b0000000000011100, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000010100, 16'b1111111111100001, 16'b1111111111111001, 16'b1111111111111100, 16'b1111111111111110, 16'b0000000000001100, 16'b1111111111111100, 16'b0000000000000001, 16'b0000000000011110, 16'b1111111111011111, 16'b1111111111101000, 16'b0000000000000001}, 
{16'b0000000000000001, 16'b1111111111111100, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111010001, 16'b1111111111011001, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111101111, 16'b0000000000000001, 16'b0000000000000000, 16'b1111111111111110, 16'b0000000000000000, 16'b1111111111111100, 16'b1111111111111100, 16'b1111111111111011, 16'b1111111111110110, 16'b0000000000010010, 16'b0000000000000000, 16'b0000000000000010, 16'b1111111111111111, 16'b1111111111111011, 16'b0000000000000000, 16'b1111111111111010, 16'b0000000000001110, 16'b1111111111011000, 16'b0000000000001110, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000001100, 16'b1111111111111111, 16'b0000000000001111}, 
{16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111101, 16'b0000000000000100, 16'b0000000000000011, 16'b1111111111101010, 16'b0000000000000000, 16'b0000000000000100, 16'b0000000000100101, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000011, 16'b0000000000010110, 16'b1111111111111101, 16'b0000000000000000, 16'b0000000000000110, 16'b1111111111111111, 16'b0000000000000001, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111101110, 16'b0000000000000010, 16'b0000000000000100, 16'b0000000000000001, 16'b1111111111111111, 16'b0000000000001101, 16'b0000000000000000, 16'b0000000000001000, 16'b1111111111100101, 16'b0000000000000110, 16'b0000000000011001, 16'b0000000000000000}, 
{16'b1111111111101001, 16'b0000000000001101, 16'b1111111111101111, 16'b0000000000000111, 16'b1111111111111001, 16'b0000000000000000, 16'b0000000000011111, 16'b1111111111110001, 16'b1111111111101101, 16'b0000000000001010, 16'b1111111111110001, 16'b1111111111111110, 16'b1111111111111111, 16'b0000000000010110, 16'b1111111111111111, 16'b1111111111101100, 16'b1111111111111111, 16'b0000000000011100, 16'b1111111111100001, 16'b1111111111111110, 16'b0000000000010100, 16'b1111111111101000, 16'b0000000000000011, 16'b1111111111111111, 16'b0000000000010001, 16'b1111111111011111, 16'b1111111111101000, 16'b1111111111110011, 16'b1111111111111111, 16'b0000000000000110, 16'b0000000000000001, 16'b0000000000001011}, 
{16'b1111111111111010, 16'b0000000000000011, 16'b1111111111111111, 16'b0000000000001001, 16'b1111111111111101, 16'b0000000000001110, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000100001, 16'b0000000000000000, 16'b0000000000001100, 16'b0000000000000000, 16'b1111111111110010, 16'b1111111111111011, 16'b1111111111111111, 16'b1111111111111110, 16'b0000000000000010, 16'b1111111111111111, 16'b1111111111110100, 16'b1111111111111111, 16'b0000000000010010, 16'b0000000000010011, 16'b1111111111111111, 16'b1111111111111110, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111001}, 
{16'b1111111111111010, 16'b0000000000000000, 16'b0000000000010001, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111000, 16'b0000000000000000, 16'b1111111111001000, 16'b0000000000001101, 16'b0000000000000000, 16'b0000000000000001, 16'b1111111111101000, 16'b0000000000000000, 16'b1111111111110111, 16'b1111111111111101, 16'b0000000000000000, 16'b0000000000000001, 16'b0000000000000000, 16'b0000000000000111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000010101, 16'b0000000000011000, 16'b1111111111110001, 16'b1111111111110110, 16'b0000000000001111, 16'b1111111111101100, 16'b0000000000000001, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000001011}, 
{16'b1111111111111000, 16'b1111111111111111, 16'b1111111111110000, 16'b1111111111110011, 16'b1111111111111111, 16'b1111111111110111, 16'b0000000000000000, 16'b0000000000000101, 16'b1111111111110000, 16'b1111111111111010, 16'b1111111111111100, 16'b0000000000000000, 16'b0000000000000001, 16'b1111111111111111, 16'b1111111111111100, 16'b0000000000000110, 16'b0000000000001110, 16'b0000000000001000, 16'b1111111111110111, 16'b0000000000000011, 16'b1111111111111111, 16'b1111111111111110, 16'b0000000000000001, 16'b0000000000000001, 16'b1111111111111011, 16'b0000000000000101, 16'b1111111111111010, 16'b0000000000000011, 16'b1111111111111111, 16'b1111111111101101, 16'b1111111111111110, 16'b0000000000001110}, 
{16'b1111111111111110, 16'b1111111111111010, 16'b0000000000000100, 16'b0000000000010000, 16'b0000000000000101, 16'b0000000000000101, 16'b0000000000000010, 16'b1111111111110011, 16'b1111111111110010, 16'b0000000000000100, 16'b0000000000000000, 16'b0000000000000010, 16'b0000000000000001, 16'b0000000000000000, 16'b0000000000001101, 16'b0000000000000000, 16'b1111111111111100, 16'b0000000000000110, 16'b1111111111111110, 16'b1111111111111101, 16'b0000000000000111, 16'b1111111111111000, 16'b1111111111111110, 16'b0000000000001000, 16'b0000000000000001, 16'b1111111111111001, 16'b1111111111110011, 16'b1111111111111111, 16'b1111111111101110, 16'b0000000000000011, 16'b0000000000000110, 16'b0000000000000000}, 
{16'b1111111111111111, 16'b1111111111111110, 16'b1111111111111111, 16'b1111111111111101, 16'b1111111111110111, 16'b1111111111110111, 16'b0000000000000100, 16'b0000000000000000, 16'b1111111111110100, 16'b0000000000001010, 16'b1111111111111110, 16'b1111111111111111, 16'b1111111111111000, 16'b0000000000000000, 16'b0000000000000001, 16'b1111111111111100, 16'b1111111111111110, 16'b1111111111111101, 16'b1111111111111010, 16'b0000000000000000, 16'b1111111111110111, 16'b0000000000000110, 16'b1111111111110010, 16'b0000000000000000, 16'b0000000000000010, 16'b0000000000000111, 16'b0000000000000001, 16'b0000000000000000, 16'b0000000000010010, 16'b0000000000000011, 16'b0000000000000000, 16'b0000000000000101}, 
{16'b1111111111111110, 16'b0000000000010000, 16'b1111111111111111, 16'b1111111111111101, 16'b1111111111110010, 16'b1111111111111011, 16'b0000000000011010, 16'b1111111111010011, 16'b1111111111101001, 16'b1111111111110011, 16'b1111111111110001, 16'b1111111111101111, 16'b1111111111111111, 16'b0000000000011110, 16'b1111111111111110, 16'b0000000000000000, 16'b1111111111110010, 16'b0000000000011100, 16'b1111111111100101, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111101010, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000011, 16'b1111111111111100, 16'b1111111111110110, 16'b1111111111111111, 16'b0000000000001011, 16'b0000000000000000, 16'b1111111111111010, 16'b0000000000000000}, 
{16'b0000000000010111, 16'b1111111111111000, 16'b0000000000001000, 16'b1111111111111101, 16'b0000000000000100, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111010, 16'b0000000000000000, 16'b0000000000000101, 16'b1111111111111111, 16'b1111111111111100, 16'b1111111111111111, 16'b0000000000001110, 16'b0000000000000001, 16'b0000000000000010, 16'b0000000000000001, 16'b1111111111111110, 16'b0000000000000001, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111101100, 16'b1111111111111111, 16'b0000000000000011, 16'b1111111111111000, 16'b1111111111110111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000100011, 16'b1111111111101101, 16'b1111111111111000}, 
{16'b1111111111111101, 16'b1111111111111001, 16'b1111111111111011, 16'b0000000000000010, 16'b0000000000001000, 16'b1111111111110111, 16'b1111111111111111, 16'b1111111111110001, 16'b0000000000000011, 16'b0000000000001000, 16'b1111111111110010, 16'b1111111111101111, 16'b0000000000000001, 16'b1111111111010100, 16'b1111111111111011, 16'b1111111111111000, 16'b1111111111110011, 16'b1111111111111111, 16'b0000000000001000, 16'b0000000000000000, 16'b1111111111111101, 16'b1111111111111101, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111100, 16'b1111111111001111, 16'b1111111111011100, 16'b1111111111101110, 16'b0000000000000011, 16'b0000000000001101, 16'b1111111111111111, 16'b0000000000001111}, 
{16'b1111111111111010, 16'b1111111111110010, 16'b0000000000001010, 16'b0000000000000100, 16'b0000000000000010, 16'b1111111111111010, 16'b1111111111111101, 16'b0000000000000110, 16'b0000000000100010, 16'b1111111111110101, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000111, 16'b1111111111111100, 16'b1111111111111110, 16'b1111111111111110, 16'b1111111111111001, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000001110, 16'b1111111111110111, 16'b1111111111111111, 16'b0000000000001000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000100001, 16'b0000000000010100, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111100101, 16'b1111111111111011, 16'b1111111111111111}, 
{16'b0000000000000000, 16'b0000000000000011, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000001110, 16'b1111111111100001, 16'b0000000000000000, 16'b1111111111111001, 16'b0000000000001011, 16'b0000000000000000, 16'b1111111111111110, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111001, 16'b0000000000010000, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111101011, 16'b0000000000000011, 16'b0000000000001011, 16'b1111111111111111, 16'b0000000000000110, 16'b1111111111111111, 16'b0000000000000100}, 
{16'b1111111111110011, 16'b0000000000000000, 16'b1111111111100001, 16'b0000000000000000, 16'b1111111111111100, 16'b1111111111111101, 16'b1111111111111111, 16'b1111111111111010, 16'b1111111111111101, 16'b1111111111111011, 16'b0000000000000011, 16'b0000000000000001, 16'b1111111111110100, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000100, 16'b1111111111111110, 16'b1111111111111110, 16'b1111111111111110, 16'b1111111111111111, 16'b0000000000010001, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000010100, 16'b0000000000001100, 16'b0000000000000010, 16'b1111111111111001, 16'b1111111111111111, 16'b0000000000000100, 16'b0000000000000011}, 
{16'b0000000000000010, 16'b0000000000000010, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111100010, 16'b0000000000000010, 16'b0000000000000001, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111110101, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111110101, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111101001, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000001000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000011101, 16'b0000000000010101, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111110001, 16'b0000000000000000, 16'b1111111111111111}, 
{16'b0000000000000100, 16'b0000000000000011, 16'b0000000000010000, 16'b1111111111110000, 16'b0000000000001000, 16'b0000000000000111, 16'b0000000000000000, 16'b0000000000001100, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000010, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000111, 16'b1111111111111111, 16'b1111111111111101, 16'b0000000000000000, 16'b0000000000000010, 16'b1111111111111100, 16'b0000000000000110, 16'b0000000000000010, 16'b1111111111011010, 16'b1111111111111000, 16'b0000000000000101, 16'b1111111111111111, 16'b1111111111011111, 16'b1111111111110111, 16'b1111111111111110, 16'b1111111111111111, 16'b1111111111111100, 16'b0000000000000000, 16'b1111111111111101}, 
{16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111010, 16'b1111111111110101, 16'b0000000000000010, 16'b0000000000000000, 16'b0000000000000110, 16'b1111111111111111, 16'b0000000000001111, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111101010, 16'b1111111111111111, 16'b0000000000001000, 16'b1111111111111111, 16'b1111111111101111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000010000, 16'b1111111111111111, 16'b1111111111100100, 16'b1111111111111111, 16'b0000000000010000, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000001000, 16'b1111111111111001, 16'b0000000000000100, 16'b0000000000000000, 16'b1111111111110011, 16'b0000000000000000, 16'b0000000000000000}, 
{16'b1111111111110010, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000011111, 16'b1111111111111000, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111101, 16'b1111111111111100, 16'b0000000000000100, 16'b0000000000001000, 16'b1111111111111101, 16'b0000000000001111, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111101101, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111010, 16'b0000000000000000, 16'b0000000000000010, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111100, 16'b1111111111110011, 16'b1111111111101101, 16'b0000000000000000, 16'b1111111111111000, 16'b0000000000000010, 16'b1111111111111111, 16'b0000000000000100}, 
{16'b1111111111100101, 16'b1111111111110101, 16'b1111111111110110, 16'b0000000000000000, 16'b0000000000100100, 16'b1111111111110001, 16'b0000000000000000, 16'b1111111111111100, 16'b1111111111100101, 16'b0000000000001000, 16'b1111111111111111, 16'b0000000000100100, 16'b0000000000000000, 16'b1111111111111100, 16'b1111111111111111, 16'b0000000000000010, 16'b1111111111111110, 16'b0000000000000000, 16'b1111111111111101, 16'b0000000000011111, 16'b0000000000000010, 16'b1111111111111101, 16'b0000000000000111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111001, 16'b1111111111111101, 16'b1111111111100010, 16'b1111111111110110, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111100}, 
{16'b0000000000001110, 16'b1111111111001100, 16'b1111111111010001, 16'b1111111111110101, 16'b0000000000101010, 16'b1111111111111111, 16'b1111111111101001, 16'b0000000000010000, 16'b0000000000000011, 16'b0000000000000000, 16'b0000000000001101, 16'b1111111111101110, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111101, 16'b0000000000000001, 16'b1111111111111001, 16'b1111111111000101, 16'b0000000000001010, 16'b0000000000010110, 16'b0000000000010000, 16'b0000000000000000, 16'b0000000000000001, 16'b1111111111100110, 16'b1111111111010111, 16'b1111111111111111, 16'b1111111111101100, 16'b1111111111100010, 16'b1111111111110011, 16'b1111111111000111, 16'b0000000000011010, 16'b0000000000011011}, 
{16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000010000, 16'b1111111111110100, 16'b0000000000000001, 16'b0000000000000100, 16'b1111111111101001, 16'b0000000000000010, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000001111, 16'b0000000000000011, 16'b0000000000000001, 16'b0000000000000011, 16'b0000000000010101, 16'b1111111111110010, 16'b0000000000000000, 16'b1111111111110101, 16'b1111111111111111, 16'b0000000000010100, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111011100, 16'b1111111111111111, 16'b1111111111110110, 16'b1111111111111100, 16'b0000000000000000, 16'b0000000000001000, 16'b0000000000000110}, 
{16'b1111111111111101, 16'b0000000000001000, 16'b1111111111101100, 16'b0000000000000001, 16'b0000000000001100, 16'b1111111111111101, 16'b1111111111111111, 16'b0000000000001010, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111011, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111101, 16'b1111111111111000, 16'b1111111111111011, 16'b1111111111111100, 16'b1111111111111011, 16'b1111111111111000, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111101, 16'b1111111111111011, 16'b0000000000011001, 16'b0000000000000000, 16'b1111111111101000, 16'b1111111111111111, 16'b0000000000000111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000010000, 16'b1111111111111111}, 
{16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111110110, 16'b1111111111001000, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111011001, 16'b0000000000000101, 16'b1111111111111001, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111101000, 16'b1111111111111101, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000010, 16'b0000000000010110, 16'b1111111111111000, 16'b1111111111101100, 16'b0000000000000000, 16'b1111111111101111, 16'b1111111111111001, 16'b1111111111110001, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111110, 16'b1111111111100001, 16'b1111111111111101, 16'b0000000000001111}, 
{16'b0000000000000111, 16'b0000000000001110, 16'b1111111111111111, 16'b0000000000001010, 16'b1111111111110010, 16'b1111111111111000, 16'b0000000000000110, 16'b0000000000000100, 16'b1111111111111100, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111101011, 16'b1111111111111111, 16'b0000000000001001, 16'b1111111111111000, 16'b0000000000000010, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000001101, 16'b1111111111101011, 16'b0000000000010001, 16'b0000000000000011, 16'b0000000000000000, 16'b0000000000001101, 16'b0000000000000000, 16'b1111111111111101, 16'b1111111111100111, 16'b1111111111111000, 16'b1111111111110101, 16'b0000000000001011}, 
{16'b0000000000000000, 16'b0000000000000000, 16'b1111111111101000, 16'b1111111111111111, 16'b0000000000001101, 16'b1111111111110110, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000001, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111110010, 16'b0000000000000110, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000010, 16'b1111111111111111, 16'b1111111111110110, 16'b0000000000000001, 16'b0000000000000000, 16'b1111111111111101, 16'b1111111111111110, 16'b0000000000010010, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111101101, 16'b1111111111101011, 16'b0000000000001111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000001, 16'b0000000000010010}, 
{16'b1111111111101010, 16'b1111111111111111, 16'b1111111111110010, 16'b0000000000000000, 16'b1111111111101001, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111011, 16'b1111111111011101, 16'b1111111111111110, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111100, 16'b1111111111110110, 16'b1111111111111001, 16'b0000000000000100, 16'b1111111111111111, 16'b1111111111111110, 16'b0000000000000000, 16'b0000000000010101, 16'b1111111111111111, 16'b0000000000001001, 16'b0000000000000101, 16'b1111111111110111, 16'b0000000000001101, 16'b1111111111111101, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000100101}, 
{16'b1111111111101011, 16'b0000000000000001, 16'b0000000000000011, 16'b1111111111111110, 16'b0000000000001111, 16'b1111111111101100, 16'b1111111111111111, 16'b0000000000010000, 16'b0000000000001010, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111011, 16'b1111111111111010, 16'b1111111111111011, 16'b1111111111111100, 16'b0000000000000101, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000001001, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000010000, 16'b0000000000000010, 16'b0000000000000000, 16'b1111111111111001, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000100}, 
{16'b1111111111111111, 16'b0000000000000000, 16'b1111111111110010, 16'b1111111111111011, 16'b0000000000010010, 16'b1111111111111111, 16'b1111111111111011, 16'b0000000000001111, 16'b1111111111111100, 16'b0000000000010010, 16'b0000000000000101, 16'b1111111111111000, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000001, 16'b1111111111111011, 16'b1111111111101111, 16'b0000000000010001, 16'b0000000000001001, 16'b0000000000101000, 16'b0000000000001100, 16'b0000000000001111, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000011, 16'b0000000000000101, 16'b1111111111100101, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111}, 
{16'b0000000000000000, 16'b1111111111111010, 16'b1111111111111001, 16'b0000000000000000, 16'b1111111111110000, 16'b0000000000000000, 16'b0000000000001100, 16'b0000000000000110, 16'b0000000000000011, 16'b1111111111111001, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111101, 16'b0000000000001100, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111101100, 16'b0000000000000000, 16'b1111111111110011, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000001, 16'b0000000000000001, 16'b0000000000001000, 16'b1111111111111011, 16'b1111111111111111, 16'b1111111111100011, 16'b0000000000000101}, 
{16'b0000000000011100, 16'b1111111111111111, 16'b0000000000000100, 16'b1111111111111001, 16'b1111111111111010, 16'b0000000000000010, 16'b0000000000001010, 16'b0000000000000000, 16'b0000000000100001, 16'b0000000000000000, 16'b1111111111111110, 16'b0000000000000001, 16'b0000000000000110, 16'b1111111111111111, 16'b0000000000000011, 16'b0000000000000110, 16'b1111111111111111, 16'b1111111111100011, 16'b1111111111111100, 16'b1111111111111111, 16'b0000000000000111, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000111, 16'b0000000000000001, 16'b1111111111101111, 16'b1111111111111001, 16'b0000000000001000, 16'b1111111111111110, 16'b0000000000010000, 16'b1111111111111111, 16'b1111111111110100}, 
{16'b0000000000000000, 16'b0000000000000110, 16'b1111111111111111, 16'b1111111111111101, 16'b1111111111101001, 16'b1111111111111111, 16'b0000000000000010, 16'b1111111111111101, 16'b0000000000001010, 16'b1111111111111101, 16'b1111111111111111, 16'b1111111111111101, 16'b1111111111111111, 16'b1111111111111101, 16'b0000000000000000, 16'b0000000000010100, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000010, 16'b0000000000001000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000010, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000001, 16'b0000000000000000, 16'b0000000000000110}, 
{16'b1111111111101100, 16'b0000000000001000, 16'b0000000000000001, 16'b1111111111111001, 16'b1111111111100110, 16'b1111111111111110, 16'b0000000000000100, 16'b1111111111100110, 16'b0000000000100000, 16'b0000000000000100, 16'b0000000000000001, 16'b0000000000000110, 16'b0000000000000010, 16'b0000000000000000, 16'b0000000000011010, 16'b1111111111111010, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111100100, 16'b0000000000000001, 16'b0000000000001001, 16'b0000000000000010, 16'b0000000000000010, 16'b1111111111010101, 16'b1111111111101010, 16'b1111111111110000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000010100, 16'b1111111111110010}, 
{16'b1111111111111111, 16'b1111111111110011, 16'b1111111111111001, 16'b1111111111100101, 16'b1111111111101111, 16'b0000000000010101, 16'b0000000000010011, 16'b1111111111110101, 16'b0000000000000010, 16'b1111111111111101, 16'b1111111111111001, 16'b1111111111101111, 16'b0000000000000110, 16'b1111111111101101, 16'b0000000000001100, 16'b1111111111111111, 16'b0000000000010101, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111110111, 16'b1111111111111101, 16'b1111111111111011, 16'b1111111111101110, 16'b0000000000000101, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111110001, 16'b0000000000010100, 16'b0000000000010001, 16'b1111111111111010, 16'b1111111111010111, 16'b0000000000001001}, 
{16'b0000000000000000, 16'b1111111111111110, 16'b1111111111111111, 16'b1111111111111001, 16'b0000000000000001, 16'b0000000000000000, 16'b0000000000000100, 16'b0000000000000000, 16'b0000000000000111, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000110, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111110111, 16'b1111111111111001, 16'b0000000000000000, 16'b0000000000001011, 16'b0000000000000011, 16'b0000000000001000, 16'b1111111111111110, 16'b1111111111110101, 16'b1111111111111111, 16'b0000000000000100, 16'b1111111111111111, 16'b0000000000000010, 16'b1111111111111111, 16'b0000000000000100, 16'b0000000000000000, 16'b0000000000000101, 16'b1111111111100111, 16'b1111111111111111}, 
{16'b0000000000010011, 16'b1111111111111111, 16'b0000000000001001, 16'b1111111111101100, 16'b1111111111110011, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000001, 16'b0000000000000000, 16'b1111111111110111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111110111, 16'b0000000000001001, 16'b1111111111111111, 16'b1111111111111110, 16'b0000000000000000, 16'b0000000000000111, 16'b1111111111110011, 16'b0000000000000111, 16'b0000000000001000, 16'b0000000000001000, 16'b1111111111111111, 16'b0000000000100011, 16'b1111111111110110, 16'b0000000000010111, 16'b1111111111111100, 16'b1111111111101000, 16'b1111111111110100, 16'b0000000000001000}, 
{16'b1111111111011101, 16'b1111111111111110, 16'b1111111111110110, 16'b1111111111111111, 16'b0000000000010000, 16'b1111111111110100, 16'b1111111111111100, 16'b0000000000001111, 16'b0000000000000110, 16'b1111111111110000, 16'b0000000000000000, 16'b1111111111111110, 16'b1111111111111111, 16'b0000000000001000, 16'b1111111111110000, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111111110, 16'b0000000000000000, 16'b1111111111110011, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111101010, 16'b0000000000000100, 16'b0000000000100111, 16'b0000000000010110, 16'b1111111111111101, 16'b1111111111110101, 16'b1111111111100011, 16'b0000000000000000, 16'b1111111111111100}, 
{16'b0000000000000001, 16'b0000000000001101, 16'b0000000000000001, 16'b1111111111110110, 16'b0000000000000000, 16'b1111111111111110, 16'b0000000000000000, 16'b0000000000001101, 16'b0000000000001101, 16'b1111111111110111, 16'b0000000000001000, 16'b0000000000000001, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111110101, 16'b0000000000010000, 16'b1111111111111101, 16'b1111111111101011, 16'b0000000000000111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000111, 16'b1111111111111011, 16'b1111111111111111, 16'b1111111111111100, 16'b0000000000000101, 16'b1111111111110111, 16'b0000000000001000, 16'b1111111111101000, 16'b0000000000000101, 16'b1111111111111111, 16'b0000000000001010}, 
{16'b1111111111111101, 16'b0000000000000000, 16'b0000000000000101, 16'b0000000000000000, 16'b1111111111111100, 16'b1111111111111111, 16'b0000000000000110, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000001, 16'b1111111111111001, 16'b0000000000000000, 16'b0000000000000111, 16'b0000000000000010, 16'b0000000000000110, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000001000, 16'b0000000000001111, 16'b1111111111111001, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111100010, 16'b1111111111111111, 16'b1111111111111011, 16'b1111111111111111, 16'b0000000000100100, 16'b0000000000000000, 16'b1111111111110010}, 
{16'b1111111111111110, 16'b1111111111111000, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000101, 16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111110, 16'b0000000000000100, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000010, 16'b0000000000010010, 16'b1111111111111001, 16'b0000000000000000, 16'b1111111111001001, 16'b1111111111111111, 16'b1111111111111100, 16'b0000000000000000, 16'b1111111111111100, 16'b0000000000000101, 16'b1111111111110001, 16'b0000000000000111, 16'b0000000000000110, 16'b1111111111111111, 16'b1111111111010010, 16'b1111111111110001, 16'b1111111111111110, 16'b1111111111111110, 16'b0000000000011000, 16'b1111111111111111, 16'b0000000000001001}, 
{16'b0000000000000011, 16'b0000000000000000, 16'b0000000000001011, 16'b1111111111111000, 16'b1111111111111011, 16'b0000000000001111, 16'b1111111111110101, 16'b0000000000000011, 16'b1111111111101100, 16'b0000000000000000, 16'b0000000000000001, 16'b1111111111111010, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111110011, 16'b0000000000011011, 16'b1111111111110000, 16'b1111111111111111, 16'b0000000000000111, 16'b1111111111111111, 16'b0000000000000100, 16'b1111111111100001, 16'b0000000000010100, 16'b1111111111111111, 16'b1111111111111000, 16'b0000000000011111, 16'b0000000000001001, 16'b1111111111110101, 16'b1111111111110111, 16'b1111111111011101, 16'b1111111111111111, 16'b0000000000000001}, 
{16'b1111111111111111, 16'b0000000000000000, 16'b1111111111111101, 16'b1111111111101110, 16'b1111111111111111, 16'b1111111111100110, 16'b0000000000000000, 16'b0000000000010011, 16'b0000000000001111, 16'b0000000000000001, 16'b0000000000000000, 16'b1111111111111000, 16'b0000000000010101, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000011011, 16'b0000000000000000, 16'b1111111111111101, 16'b1111111111111100, 16'b1111111111101011, 16'b0000000000001000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000010, 16'b1111111111111011, 16'b1111111111100010, 16'b0000000000010001, 16'b1111111111100011, 16'b0000000000000011, 16'b1111111111111010, 16'b0000000000000000}, 
{16'b0000000000000011, 16'b0000000000001011, 16'b0000000000000000, 16'b1111111111111111, 16'b1111111111100010, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000001111, 16'b0000000000010001, 16'b1111111111111111, 16'b1111111111111111, 16'b1111111111111111, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b1111111111111111, 16'b0000000000001010, 16'b1111111111111001, 16'b1111111111100100, 16'b1111111111111101, 16'b1111111111111001, 16'b1111111111111001, 16'b1111111111111011, 16'b1111111111111111, 16'b1111111111111011, 16'b1111111111111110, 16'b1111111111111111, 16'b0000000000001001, 16'b1111111111111111, 16'b0000000000011101}
};

localparam logic signed [15:0] bias [32] = '{
16'b0000000001011110,  // 1.474280834197998
16'b0000000000101100,  // 0.6914801001548767
16'b0000000001011100,  // 1.4406442642211914
16'b0000000001011010,  // 1.408045768737793
16'b0000000000111111,  // 0.9864811301231384
16'b0000000000110111,  // 0.8636202812194824
16'b1111111111011000,  // -0.6153604388237
16'b0000000000011110,  // 0.4839226007461548
16'b0000000000011111,  // 0.4862793982028961
16'b0000000000010111,  // 0.37162142992019653
16'b0000000000011101,  // 0.45989668369293213
16'b0000000001010011,  // 1.2998151779174805
16'b1111111110111110,  // -1.016528844833374
16'b1111111111101001,  // -0.35249894857406616
16'b0000000000011100,  // 0.44582197070121765
16'b1111111111111000,  // -0.1119980737566948
16'b1111111111111011,  // -0.06717441976070404
16'b0000000000000000,  // 0.00487547367811203
16'b0000000000001100,  // 0.1946917623281479
16'b1111111111001110,  // -0.7796769738197327
16'b0000000000101110,  // 0.7287401556968689
16'b0000000001101101,  // 1.714877724647522
16'b1111111110011001,  // -1.5971007347106934
16'b0000000000000100,  // 0.07393483817577362
16'b0000000000010100,  // 0.3225609362125397
16'b0000000000110110,  // 0.8453295230865479
16'b0000000000111001,  // 0.898597240447998
16'b0000000000010000,  // 0.2548799514770508
16'b0000000000111110,  // 0.9735668301582336
16'b0000000001001000,  // 1.1261906623840332
16'b0000000000011100,  // 0.44768181443214417
16'b1111111101101000   // -2.3676068782806396
};
endpackage