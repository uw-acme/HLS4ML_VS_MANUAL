// Width: 6
// NFRAC: 3
package dense_3_6_3;

localparam logic signed [5:0] weights [32][32] = '{ 
{6'b111111, 6'b111100, 6'b111100, 6'b111110, 6'b000010, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b000001, 6'b111011, 6'b111111, 6'b000110, 6'b111110, 6'b111000, 6'b111111, 6'b000000, 6'b000011, 6'b111101, 6'b110111, 6'b111111, 6'b000000, 6'b111100, 6'b000000, 6'b001000, 6'b110100, 6'b111110, 6'b111100, 6'b111110, 6'b000011, 6'b111110}, 
{6'b000101, 6'b001101, 6'b000011, 6'b111010, 6'b000001, 6'b111101, 6'b111111, 6'b001000, 6'b000000, 6'b111111, 6'b111111, 6'b111011, 6'b111110, 6'b000100, 6'b101111, 6'b111100, 6'b111111, 6'b111111, 6'b111111, 6'b111110, 6'b111101, 6'b111101, 6'b000000, 6'b111111, 6'b111111, 6'b110111, 6'b000000, 6'b000011, 6'b111111, 6'b111010, 6'b000000, 6'b000000}, 
{6'b111000, 6'b000001, 6'b000000, 6'b000010, 6'b111010, 6'b000000, 6'b000000, 6'b111001, 6'b000100, 6'b111101, 6'b111101, 6'b110100, 6'b111101, 6'b000100, 6'b000010, 6'b111111, 6'b111111, 6'b111111, 6'b111001, 6'b000000, 6'b000000, 6'b000000, 6'b000001, 6'b000111, 6'b000000, 6'b111001, 6'b000110, 6'b000000, 6'b000001, 6'b111111, 6'b000000, 6'b010010}, 
{6'b000110, 6'b111111, 6'b111110, 6'b001010, 6'b001001, 6'b000000, 6'b000000, 6'b000110, 6'b111100, 6'b111111, 6'b111001, 6'b000000, 6'b000010, 6'b111010, 6'b000000, 6'b111110, 6'b111111, 6'b111101, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b001001, 6'b000101, 6'b000101, 6'b000011, 6'b000101, 6'b000000, 6'b111111, 6'b000111, 6'b000011, 6'b111110}, 
{6'b001000, 6'b111111, 6'b111010, 6'b110011, 6'b000111, 6'b000000, 6'b111001, 6'b111011, 6'b111111, 6'b110011, 6'b101110, 6'b000111, 6'b001010, 6'b001000, 6'b110110, 6'b110011, 6'b000000, 6'b111101, 6'b000011, 6'b000010, 6'b111100, 6'b111111, 6'b001011, 6'b101010, 6'b000001, 6'b110101, 6'b000001, 6'b111100, 6'b111011, 6'b111111, 6'b000001, 6'b001001}, 
{6'b000000, 6'b111111, 6'b111011, 6'b111011, 6'b000101, 6'b000000, 6'b111011, 6'b111101, 6'b111001, 6'b111110, 6'b111111, 6'b000010, 6'b000000, 6'b000101, 6'b110111, 6'b111101, 6'b000001, 6'b111011, 6'b111100, 6'b111111, 6'b000000, 6'b000100, 6'b000111, 6'b111111, 6'b111111, 6'b000110, 6'b110111, 6'b111111, 6'b111100, 6'b111111, 6'b111111, 6'b000000}, 
{6'b000001, 6'b111010, 6'b000001, 6'b111111, 6'b111111, 6'b000010, 6'b111110, 6'b110101, 6'b111111, 6'b111100, 6'b111000, 6'b000111, 6'b000000, 6'b001010, 6'b001101, 6'b000000, 6'b111111, 6'b111010, 6'b111111, 6'b000100, 6'b110011, 6'b000010, 6'b000101, 6'b000000, 6'b000010, 6'b010011, 6'b111001, 6'b111110, 6'b111100, 6'b000111, 6'b111111, 6'b111101}, 
{6'b110110, 6'b000000, 6'b110101, 6'b000110, 6'b010000, 6'b000001, 6'b000000, 6'b000000, 6'b111111, 6'b000010, 6'b010100, 6'b111111, 6'b000110, 6'b001001, 6'b001100, 6'b010000, 6'b000000, 6'b111000, 6'b000101, 6'b111111, 6'b110101, 6'b111100, 6'b000000, 6'b111110, 6'b110111, 6'b011110, 6'b111100, 6'b000000, 6'b000000, 6'b001110, 6'b000001, 6'b000110}, 
{6'b000110, 6'b111111, 6'b000000, 6'b111111, 6'b000001, 6'b111111, 6'b111111, 6'b000010, 6'b000011, 6'b111011, 6'b000010, 6'b000010, 6'b000000, 6'b000101, 6'b111100, 6'b110011, 6'b000000, 6'b111111, 6'b111111, 6'b111000, 6'b111111, 6'b000000, 6'b111100, 6'b111111, 6'b111110, 6'b000010, 6'b000101, 6'b111110, 6'b111111, 6'b111111, 6'b000000, 6'b111001}, 
{6'b111101, 6'b000110, 6'b000000, 6'b000000, 6'b001100, 6'b000101, 6'b111111, 6'b110111, 6'b000001, 6'b110100, 6'b101001, 6'b111111, 6'b000000, 6'b000110, 6'b000001, 6'b000000, 6'b111010, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b111111, 6'b111010, 6'b000000, 6'b111111, 6'b010001, 6'b000101, 6'b111111, 6'b111110, 6'b001010, 6'b111111, 6'b111110}, 
{6'b110111, 6'b000010, 6'b111111, 6'b111111, 6'b111100, 6'b111001, 6'b000000, 6'b000010, 6'b111111, 6'b111101, 6'b110110, 6'b000011, 6'b000100, 6'b000000, 6'b001101, 6'b110111, 6'b000001, 6'b111001, 6'b000100, 6'b111111, 6'b111111, 6'b000001, 6'b000001, 6'b000000, 6'b111000, 6'b000000, 6'b110111, 6'b111111, 6'b111111, 6'b001010, 6'b111100, 6'b000000}, 
{6'b111111, 6'b000001, 6'b000000, 6'b000110, 6'b111110, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b001010, 6'b001011, 6'b000000, 6'b111010, 6'b110100, 6'b111111, 6'b000000, 6'b000000, 6'b111110, 6'b111000, 6'b000110, 6'b000000, 6'b000101, 6'b111111, 6'b001000, 6'b000001, 6'b000100, 6'b000111, 6'b111111, 6'b111001, 6'b111000, 6'b111111, 6'b110101}, 
{6'b111100, 6'b111111, 6'b000001, 6'b111001, 6'b000001, 6'b111111, 6'b111100, 6'b111111, 6'b111101, 6'b000000, 6'b000001, 6'b111110, 6'b000000, 6'b000011, 6'b110101, 6'b111100, 6'b000011, 6'b111101, 6'b000000, 6'b111111, 6'b000011, 6'b000000, 6'b111111, 6'b000000, 6'b000100, 6'b111110, 6'b000000, 6'b111000, 6'b111100, 6'b111111, 6'b000010, 6'b000000}, 
{6'b110111, 6'b000110, 6'b111111, 6'b111111, 6'b111111, 6'b000010, 6'b111111, 6'b001100, 6'b111111, 6'b111111, 6'b000011, 6'b000000, 6'b000000, 6'b000000, 6'b000001, 6'b000101, 6'b000010, 6'b000010, 6'b111111, 6'b000100, 6'b000001, 6'b000000, 6'b111111, 6'b000100, 6'b111110, 6'b111010, 6'b111110, 6'b111111, 6'b000001, 6'b000000, 6'b000011, 6'b000111}, 
{6'b111111, 6'b111001, 6'b000000, 6'b111111, 6'b001110, 6'b111100, 6'b110110, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b000110, 6'b000101, 6'b000000, 6'b000000, 6'b111101, 6'b000000, 6'b111111, 6'b000000, 6'b000001, 6'b111111, 6'b000000, 6'b000100, 6'b000000, 6'b111111, 6'b111001, 6'b000011, 6'b111111, 6'b111111, 6'b111110, 6'b111111, 6'b111110}, 
{6'b000000, 6'b111110, 6'b111101, 6'b111100, 6'b110111, 6'b001001, 6'b000000, 6'b000010, 6'b000100, 6'b000000, 6'b111111, 6'b000111, 6'b000011, 6'b111010, 6'b111101, 6'b111111, 6'b111001, 6'b111111, 6'b000000, 6'b111111, 6'b000010, 6'b111101, 6'b000000, 6'b000001, 6'b111111, 6'b111010, 6'b000010, 6'b000000, 6'b000000, 6'b000000, 6'b111010, 6'b000000}, 
{6'b111100, 6'b111101, 6'b000001, 6'b111110, 6'b111110, 6'b000001, 6'b111111, 6'b000000, 6'b000010, 6'b111111, 6'b000001, 6'b111101, 6'b111111, 6'b111111, 6'b000001, 6'b111111, 6'b000111, 6'b111111, 6'b000011, 6'b111101, 6'b000010, 6'b000001, 6'b000001, 6'b000000, 6'b111110, 6'b111011, 6'b111011, 6'b000001, 6'b111110, 6'b000000, 6'b111111, 6'b000011}, 
{6'b111111, 6'b111001, 6'b111001, 6'b111111, 6'b001010, 6'b111110, 6'b000000, 6'b000111, 6'b111101, 6'b000000, 6'b111001, 6'b111000, 6'b000111, 6'b000010, 6'b111110, 6'b111011, 6'b000010, 6'b000000, 6'b111100, 6'b000000, 6'b000001, 6'b111110, 6'b000100, 6'b110000, 6'b000000, 6'b000011, 6'b111111, 6'b000000, 6'b111100, 6'b111111, 6'b111100, 6'b111111}, 
{6'b000011, 6'b000101, 6'b001000, 6'b111100, 6'b000110, 6'b000100, 6'b000000, 6'b000111, 6'b000101, 6'b111110, 6'b001011, 6'b111010, 6'b001001, 6'b000111, 6'b101110, 6'b111111, 6'b000000, 6'b000000, 6'b000100, 6'b110111, 6'b000011, 6'b111100, 6'b111000, 6'b111101, 6'b000101, 6'b110101, 6'b111010, 6'b111111, 6'b111111, 6'b110110, 6'b000110, 6'b000000}, 
{6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b111010, 6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b000010, 6'b111111, 6'b000001, 6'b111010, 6'b000001, 6'b111111, 6'b000010, 6'b000111, 6'b111010, 6'b000000, 6'b111110, 6'b000010, 6'b000011, 6'b111110, 6'b111011, 6'b000000, 6'b001101, 6'b111111, 6'b111111, 6'b000101, 6'b000000, 6'b001101}, 
{6'b110111, 6'b000000, 6'b111100, 6'b000110, 6'b000001, 6'b111111, 6'b111111, 6'b111111, 6'b111011, 6'b111111, 6'b000000, 6'b110111, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b111110, 6'b000000, 6'b000000, 6'b000010, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b001001, 6'b111111, 6'b111111, 6'b111111, 6'b000010, 6'b111111}, 
{6'b111111, 6'b111101, 6'b000011, 6'b000000, 6'b111010, 6'b000000, 6'b000100, 6'b111111, 6'b000000, 6'b111110, 6'b000001, 6'b000000, 6'b000101, 6'b110111, 6'b111110, 6'b111111, 6'b000011, 6'b111001, 6'b000000, 6'b110011, 6'b111111, 6'b111110, 6'b111111, 6'b000100, 6'b111110, 6'b111011, 6'b000001, 6'b000000, 6'b000110, 6'b001000, 6'b111010, 6'b111000}, 
{6'b000001, 6'b000000, 6'b111001, 6'b111111, 6'b111111, 6'b000000, 6'b000001, 6'b000110, 6'b000000, 6'b000000, 6'b000001, 6'b110111, 6'b111110, 6'b110110, 6'b000111, 6'b000000, 6'b111111, 6'b110101, 6'b111111, 6'b111110, 6'b111111, 6'b000000, 6'b000000, 6'b111101, 6'b000000, 6'b000110, 6'b000110, 6'b000110, 6'b000100, 6'b000000, 6'b000001, 6'b001100}, 
{6'b111111, 6'b111100, 6'b000110, 6'b111110, 6'b000001, 6'b000010, 6'b111111, 6'b111011, 6'b111110, 6'b110110, 6'b000111, 6'b000000, 6'b000110, 6'b001010, 6'b111110, 6'b110010, 6'b111110, 6'b000111, 6'b111011, 6'b111100, 6'b000000, 6'b000000, 6'b110111, 6'b111100, 6'b111111, 6'b111110, 6'b000001, 6'b001011, 6'b000011, 6'b111111, 6'b000001, 6'b000000}, 
{6'b000000, 6'b000111, 6'b000000, 6'b000100, 6'b001101, 6'b111101, 6'b111111, 6'b111111, 6'b000100, 6'b111100, 6'b111111, 6'b000101, 6'b000000, 6'b000000, 6'b100111, 6'b111110, 6'b000000, 6'b000011, 6'b111111, 6'b000100, 6'b111111, 6'b111101, 6'b110111, 6'b000010, 6'b000100, 6'b101110, 6'b111111, 6'b000000, 6'b001000, 6'b110011, 6'b000000, 6'b111111}, 
{6'b000000, 6'b111010, 6'b000000, 6'b111111, 6'b000000, 6'b001000, 6'b110100, 6'b000000, 6'b000110, 6'b111010, 6'b111111, 6'b000000, 6'b111111, 6'b000010, 6'b000001, 6'b111111, 6'b000001, 6'b000000, 6'b000000, 6'b000110, 6'b111111, 6'b111000, 6'b110110, 6'b111100, 6'b110110, 6'b000011, 6'b001001, 6'b000101, 6'b111111, 6'b111010, 6'b111011, 6'b000000}, 
{6'b000000, 6'b111000, 6'b111111, 6'b000010, 6'b111000, 6'b000010, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b000100, 6'b111111, 6'b000000, 6'b000000, 6'b000010, 6'b111111, 6'b000000, 6'b111111, 6'b111010, 6'b110111, 6'b111111, 6'b110111, 6'b111011, 6'b111010, 6'b001110, 6'b000000, 6'b111111, 6'b000101, 6'b001110, 6'b000110, 6'b101111, 6'b111101}, 
{6'b000110, 6'b111111, 6'b000100, 6'b111111, 6'b000111, 6'b111101, 6'b000001, 6'b000110, 6'b000100, 6'b110111, 6'b111111, 6'b000001, 6'b000001, 6'b111111, 6'b000001, 6'b000000, 6'b000101, 6'b000000, 6'b000101, 6'b111110, 6'b111101, 6'b111110, 6'b111111, 6'b000100, 6'b111100, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b000100, 6'b111010, 6'b111111}, 
{6'b111111, 6'b111111, 6'b111000, 6'b000100, 6'b000011, 6'b111110, 6'b111111, 6'b111100, 6'b000000, 6'b111111, 6'b111011, 6'b111100, 6'b000111, 6'b000000, 6'b111101, 6'b111111, 6'b000011, 6'b111111, 6'b111111, 6'b111100, 6'b000101, 6'b000000, 6'b000010, 6'b111111, 6'b000010, 6'b000000, 6'b000000, 6'b000011, 6'b111100, 6'b111111, 6'b000010, 6'b111110}, 
{6'b111111, 6'b111011, 6'b001001, 6'b111110, 6'b000011, 6'b111011, 6'b000000, 6'b000000, 6'b111000, 6'b111111, 6'b111110, 6'b000000, 6'b111010, 6'b000010, 6'b000011, 6'b000001, 6'b000001, 6'b111111, 6'b110100, 6'b111111, 6'b111111, 6'b000010, 6'b111110, 6'b111111, 6'b000011, 6'b111111, 6'b111111, 6'b000110, 6'b111001, 6'b111011, 6'b000101, 6'b000000}, 
{6'b000110, 6'b000011, 6'b000000, 6'b111101, 6'b111110, 6'b111111, 6'b000000, 6'b111110, 6'b111110, 6'b111110, 6'b000000, 6'b000010, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b111101, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b000001, 6'b000000, 6'b000000, 6'b110110, 6'b111100, 6'b000000, 6'b000000, 6'b000000, 6'b111101, 6'b000000}, 
{6'b000011, 6'b101111, 6'b111111, 6'b111110, 6'b111100, 6'b111111, 6'b000000, 6'b001000, 6'b111111, 6'b111111, 6'b000001, 6'b110101, 6'b000000, 6'b111000, 6'b001011, 6'b111111, 6'b111100, 6'b110111, 6'b111111, 6'b110100, 6'b110011, 6'b111111, 6'b000000, 6'b000000, 6'b000011, 6'b111111, 6'b111011, 6'b111110, 6'b111111, 6'b000000, 6'b111111, 6'b110100}
};

localparam logic signed [5:0] bias [32] = '{
6'b000100,  // 0.5280959606170654
6'b000110,  // 0.8414360880851746
6'b000011,  // 0.397830605506897
6'b000011,  // 0.4105983078479767
6'b100010,  // -3.657735586166382
6'b111000,  // -0.8977976441383362
6'b001101,  // 1.7051936388015747
6'b110101,  // -1.2765135765075684
6'b111011,  // -0.5837795734405518
6'b010101,  // 2.699671983718872
6'b000001,  // 0.2170683741569519
6'b000111,  // 0.8814588785171509
6'b101010,  // -2.634300947189331
6'b110000,  // -1.877297282218933
6'b001101,  // 1.6625694036483765
6'b010101,  // 2.7459704875946045
6'b111100,  // -0.47838035225868225
6'b001101,  // 1.6984987258911133
6'b000110,  // 0.8548859357833862
6'b001000,  // 1.0045719146728516
6'b001011,  // 1.4197649955749512
6'b000110,  // 0.832463800907135
6'b000100,  // 0.5434179306030273
6'b000111,  // 0.9277304410934448
6'b111101,  // -0.3426123857498169
6'b111011,  // -0.5587119460105896
6'b111011,  // -0.6208624839782715
6'b110101,  // -1.2802538871765137
6'b000000,  // 0.05940237268805504
6'b111001,  // -0.8213341236114502
6'b000111,  // 0.8783953189849854
6'b111000   // -0.949700653553009
};
endpackage