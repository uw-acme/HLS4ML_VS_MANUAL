// Width: 10
// NFRAC: 5
package dense_1_10_5;

localparam logic signed [9:0] weights [16][64] = '{ 
{10'b0000001000, 10'b1111101011, 10'b1111111010, 10'b1111111000, 10'b1111110011, 10'b0000000011, 10'b1111011110, 10'b0000000000, 10'b0000000001, 10'b0000001000, 10'b0000000000, 10'b1111110011, 10'b1111111111, 10'b0000000110, 10'b0000000001, 10'b1111110111, 10'b0000000111, 10'b0000000001, 10'b0000000000, 10'b1111111111, 10'b0000001100, 10'b1111110101, 10'b1111111111, 10'b0000001111, 10'b1111110101, 10'b1111101010, 10'b1111110111, 10'b1111111001, 10'b1111111100, 10'b1111111111, 10'b0000000001, 10'b0000000111, 10'b0000000110, 10'b1111111111, 10'b0000000000, 10'b0000001001, 10'b1111111111, 10'b1111110111, 10'b0000000000, 10'b0000000110, 10'b1111111111, 10'b0000001000, 10'b1111110111, 10'b0000011101, 10'b1111111111, 10'b0000001110, 10'b0000000000, 10'b0000000101, 10'b0000000110, 10'b1111111111, 10'b0000000000, 10'b0000000101, 10'b0000000110, 10'b0000000010, 10'b1111111100, 10'b1111110110, 10'b0000010001, 10'b1111110000, 10'b0000001110, 10'b1111110100, 10'b0000011001, 10'b1111111111, 10'b0000000000, 10'b0000000010}, 
{10'b0000000000, 10'b1111110101, 10'b1111111011, 10'b1111110111, 10'b1111110101, 10'b0000000011, 10'b1111100111, 10'b1111111111, 10'b1111111000, 10'b0000000101, 10'b0000000000, 10'b1111111101, 10'b0000000110, 10'b0000000000, 10'b1111111111, 10'b0000000110, 10'b1111111111, 10'b0000000000, 10'b1111111010, 10'b1111110111, 10'b0000001110, 10'b1111111101, 10'b0000000001, 10'b0000010110, 10'b0000001000, 10'b1111111000, 10'b1111111000, 10'b1111111111, 10'b1111111100, 10'b1111110011, 10'b1111111110, 10'b0000001110, 10'b0000001000, 10'b0000010001, 10'b0000010100, 10'b0000000001, 10'b1111111100, 10'b1111110010, 10'b0000000001, 10'b0000000110, 10'b0000000000, 10'b0000000110, 10'b1111111001, 10'b0000001000, 10'b0000000101, 10'b0000000001, 10'b1111110101, 10'b0000000010, 10'b0000001000, 10'b0000000000, 10'b0000000000, 10'b0000100101, 10'b1111111101, 10'b1111111100, 10'b1111111110, 10'b1111111111, 10'b0000001000, 10'b1111110100, 10'b0000011111, 10'b0000000000, 10'b0000010000, 10'b0000000111, 10'b0000011010, 10'b0000000100}, 
{10'b1111111111, 10'b0000000000, 10'b1111111101, 10'b1111111010, 10'b1111111010, 10'b0000000001, 10'b0000101111, 10'b1111111111, 10'b1111010111, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b1111111000, 10'b0000000000, 10'b1111111111, 10'b0000000101, 10'b0000011100, 10'b1111111111, 10'b0000000010, 10'b0000000000, 10'b0000001101, 10'b1111101000, 10'b0000010010, 10'b1111101001, 10'b0000011110, 10'b1111110100, 10'b1111111000, 10'b1111101001, 10'b0000101000, 10'b0000001000, 10'b0000000000, 10'b0000010000, 10'b0000100000, 10'b1111011001, 10'b1111111100, 10'b0000000001, 10'b1111111000, 10'b0000011100, 10'b1111111110, 10'b0000001010, 10'b0000001010, 10'b0000001011, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b0000000101, 10'b1111110111, 10'b1111111010, 10'b1111111111, 10'b0000001100, 10'b1111111010, 10'b0000000100, 10'b1111111111, 10'b0000000100, 10'b1111111010, 10'b1111111111, 10'b1111110110, 10'b1111101010, 10'b1111111111, 10'b0000000000, 10'b0000110001, 10'b0000000000, 10'b1111111111, 10'b1111110110}, 
{10'b1111110001, 10'b1111110100, 10'b1111101001, 10'b0000001001, 10'b1111110101, 10'b1111010100, 10'b1111111100, 10'b1111110110, 10'b0000000111, 10'b1111111111, 10'b0000101000, 10'b1111111100, 10'b1111100110, 10'b0000010010, 10'b0000000000, 10'b1111111111, 10'b1111110001, 10'b1111111111, 10'b0000000000, 10'b1111111000, 10'b1111011011, 10'b1111111100, 10'b1111101001, 10'b0000000110, 10'b1111110011, 10'b1111100010, 10'b0000001010, 10'b0000010111, 10'b0000101001, 10'b1111110001, 10'b1111101101, 10'b0000000010, 10'b0000010000, 10'b1111100101, 10'b1111110101, 10'b0000000000, 10'b1111101000, 10'b0000000111, 10'b1111110001, 10'b0000000011, 10'b0000001110, 10'b0000000101, 10'b0000000000, 10'b0000000000, 10'b0000010001, 10'b1111111001, 10'b1111111111, 10'b1111110100, 10'b1111111111, 10'b1111111100, 10'b1111101100, 10'b0000000010, 10'b1111111111, 10'b0000000110, 10'b0000001010, 10'b0000010100, 10'b1111100001, 10'b1111100010, 10'b1111101001, 10'b0000011011, 10'b0000110111, 10'b1111100011, 10'b1111111110, 10'b0000001101}, 
{10'b0000001010, 10'b1111101100, 10'b1111110111, 10'b1111111111, 10'b1111111011, 10'b0000001010, 10'b0000000110, 10'b1111111111, 10'b1111101100, 10'b1111111000, 10'b1111110100, 10'b0000000001, 10'b0000000000, 10'b0000000000, 10'b1111111110, 10'b0000001011, 10'b0000000100, 10'b1111110011, 10'b0000000000, 10'b0000000000, 10'b0000000110, 10'b1111111100, 10'b0000000010, 10'b1111111111, 10'b0000100010, 10'b1111111010, 10'b1111110111, 10'b1111110011, 10'b0000000000, 10'b0000000101, 10'b0000000011, 10'b0000001000, 10'b1111111111, 10'b0000000010, 10'b0000000100, 10'b1111111111, 10'b0000000000, 10'b0000011100, 10'b1111110110, 10'b1111111101, 10'b0000001101, 10'b0000000111, 10'b1111110000, 10'b0000000000, 10'b1111011101, 10'b1111111111, 10'b1111111100, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b0000000110, 10'b1111111111, 10'b0000001010, 10'b1111111001, 10'b1111101000, 10'b1111110001, 10'b1111101111, 10'b1111101100, 10'b0000010111, 10'b0000101011, 10'b0000011001, 10'b0000000011, 10'b1111111111}, 
{10'b1111110001, 10'b1111101011, 10'b0000000000, 10'b0000001001, 10'b0000001001, 10'b1111111001, 10'b0000010010, 10'b1111111111, 10'b0000000111, 10'b1111111111, 10'b1111111111, 10'b1111111101, 10'b1111111010, 10'b0000010010, 10'b1111111101, 10'b0000000000, 10'b1111101100, 10'b1111110100, 10'b0000000000, 10'b1111111111, 10'b1111111110, 10'b1111110101, 10'b1111110101, 10'b0000001110, 10'b1111110101, 10'b1111111111, 10'b0000001000, 10'b1111111101, 10'b1111100010, 10'b1111111111, 10'b1111111101, 10'b1111111111, 10'b1111111111, 10'b0000000001, 10'b0000000100, 10'b0000001011, 10'b0000000000, 10'b1111111100, 10'b1111110111, 10'b1111111111, 10'b1111111010, 10'b1111101111, 10'b0000001100, 10'b0000000000, 10'b0000010011, 10'b0000000000, 10'b1111111111, 10'b0000000011, 10'b1111110010, 10'b0000000111, 10'b0000000000, 10'b1111111100, 10'b1111110100, 10'b0000001100, 10'b1111111111, 10'b0000001011, 10'b0000000110, 10'b0000000110, 10'b1111111111, 10'b1111111111, 10'b1111100110, 10'b1111111011, 10'b1111111110, 10'b1111111111}, 
{10'b1111110110, 10'b1111110101, 10'b1111110010, 10'b1111111101, 10'b1111111011, 10'b0000000011, 10'b1111101001, 10'b1111111011, 10'b1111111000, 10'b1111111111, 10'b1111110110, 10'b0000001011, 10'b0000000001, 10'b0000000100, 10'b0000001001, 10'b0000000000, 10'b0000011001, 10'b0000000010, 10'b0000000111, 10'b0000001000, 10'b1111111010, 10'b0000001011, 10'b1111111000, 10'b1111101111, 10'b0000000101, 10'b0000010000, 10'b1111111111, 10'b0000000001, 10'b1111100001, 10'b0000001001, 10'b0000001000, 10'b1111110100, 10'b0000001111, 10'b0000010101, 10'b0000000000, 10'b0000001010, 10'b1111111111, 10'b0000001001, 10'b0000000110, 10'b0000000000, 10'b1111111100, 10'b1111110100, 10'b0000000100, 10'b0000001111, 10'b0000010000, 10'b1111111010, 10'b1111111101, 10'b1111111001, 10'b1111111011, 10'b0000000011, 10'b0000000000, 10'b0000000001, 10'b0000000000, 10'b0000000101, 10'b1111111010, 10'b0000011000, 10'b0000001011, 10'b1111111111, 10'b0000001100, 10'b0000000110, 10'b1111001011, 10'b1111101101, 10'b1111111010, 10'b1111111111}, 
{10'b0000000000, 10'b0000000111, 10'b1111111111, 10'b1111111111, 10'b1111110101, 10'b1111111111, 10'b1111110111, 10'b0000000000, 10'b0000000000, 10'b0000001100, 10'b0000000000, 10'b1111110011, 10'b1111111101, 10'b0000000000, 10'b1111111110, 10'b1111110001, 10'b1111100100, 10'b1111111111, 10'b1111101100, 10'b1111110001, 10'b1111110011, 10'b0000001011, 10'b0000000001, 10'b1111111011, 10'b1111110010, 10'b0000000100, 10'b0000000000, 10'b0000001111, 10'b0000011001, 10'b1111111110, 10'b0000000000, 10'b0000000111, 10'b1111101010, 10'b1111110100, 10'b0000000001, 10'b0000000010, 10'b1111110111, 10'b0000000111, 10'b0000000100, 10'b1111111011, 10'b1111110010, 10'b1111111110, 10'b0000000001, 10'b1111111010, 10'b0000000001, 10'b0000000111, 10'b1111111100, 10'b0000000000, 10'b0000000000, 10'b1111111001, 10'b1111110011, 10'b0000001101, 10'b0000000100, 10'b1111111010, 10'b0000000100, 10'b1111111110, 10'b1111110000, 10'b1111111011, 10'b1111111110, 10'b1111111101, 10'b0000011010, 10'b0000000110, 10'b1111111110, 10'b1111111111}, 
{10'b0000000000, 10'b0000010010, 10'b1111101101, 10'b1111111000, 10'b0000001010, 10'b1111111001, 10'b0000100110, 10'b1111110110, 10'b1111111111, 10'b0000001001, 10'b0000001000, 10'b1111111111, 10'b1111111110, 10'b1111110000, 10'b0000001001, 10'b0000000101, 10'b1111111001, 10'b1111111111, 10'b0000000000, 10'b0000000000, 10'b0000001000, 10'b1111110001, 10'b0000001100, 10'b0000010011, 10'b1111111101, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b0000010111, 10'b0000000000, 10'b1111110111, 10'b0000000000, 10'b0000001100, 10'b1111100110, 10'b1111101110, 10'b0000000110, 10'b0000000100, 10'b1111101101, 10'b1111111001, 10'b1111111001, 10'b0000001100, 10'b0000001100, 10'b0000000000, 10'b1111110111, 10'b0000000000, 10'b0000001100, 10'b1111111110, 10'b1111111111, 10'b0000000000, 10'b0000000111, 10'b1111111110, 10'b1111111001, 10'b0000001011, 10'b1111111001, 10'b0000001000, 10'b0000010010, 10'b0000000001, 10'b0000001000, 10'b1111110011, 10'b1111110100, 10'b0000011010, 10'b1111111011, 10'b0000000001, 10'b1111111101}, 
{10'b0000000000, 10'b1111110001, 10'b0000001011, 10'b1111110110, 10'b1111111111, 10'b0000000110, 10'b1111101101, 10'b0000000110, 10'b0000001111, 10'b0000000100, 10'b0000001011, 10'b0000001010, 10'b1111110110, 10'b1111111101, 10'b1111111110, 10'b0000000000, 10'b1111100001, 10'b0000001010, 10'b1111111110, 10'b0000000000, 10'b1111110100, 10'b0000000010, 10'b0000000100, 10'b1111111111, 10'b1111110001, 10'b1111111110, 10'b1111111101, 10'b0000100111, 10'b1111101010, 10'b0000000010, 10'b0000000011, 10'b1111111110, 10'b1111111000, 10'b0000000011, 10'b1111111101, 10'b1111111011, 10'b1111111010, 10'b1111111001, 10'b1111111111, 10'b1111110110, 10'b0000001010, 10'b0000000011, 10'b0000001111, 10'b0000000010, 10'b0000000001, 10'b1111110110, 10'b0000000000, 10'b1111111111, 10'b1111111111, 10'b0000000110, 10'b0000000101, 10'b0000001001, 10'b1111111111, 10'b1111110110, 10'b0000000000, 10'b0000000000, 10'b0000001010, 10'b1111111001, 10'b1111101110, 10'b0000010001, 10'b1111110110, 10'b0000100101, 10'b1111111111, 10'b1111110100}, 
{10'b1111101101, 10'b1111111111, 10'b1111110010, 10'b0000000111, 10'b0000001000, 10'b1111111100, 10'b0000010000, 10'b1111111010, 10'b1111110000, 10'b1111110100, 10'b1111110111, 10'b1111110000, 10'b1111111000, 10'b0000000110, 10'b0000000000, 10'b0000000000, 10'b0000011010, 10'b1111111110, 10'b1111111111, 10'b0000001101, 10'b0000001001, 10'b1111101101, 10'b1111110011, 10'b0000000110, 10'b1111110010, 10'b1111111111, 10'b1111110111, 10'b1111110101, 10'b1111110010, 10'b0000001001, 10'b0000000111, 10'b1111111011, 10'b1111111101, 10'b1111100000, 10'b1111111010, 10'b0000000001, 10'b1111111011, 10'b1111110110, 10'b1111111111, 10'b0000000011, 10'b1111111100, 10'b1111111111, 10'b1111111110, 10'b1111101010, 10'b0000000000, 10'b0000000000, 10'b0000001010, 10'b1111111100, 10'b0000001101, 10'b1111111001, 10'b0000001001, 10'b1111111111, 10'b0000000111, 10'b1111110011, 10'b1111111111, 10'b0000010000, 10'b0000001010, 10'b0000001001, 10'b0000000000, 10'b1111110011, 10'b1111110110, 10'b1111101010, 10'b1111111111, 10'b0000000011}, 
{10'b0000001001, 10'b0000000000, 10'b0000000100, 10'b1111111111, 10'b0000000100, 10'b1111111011, 10'b0000000111, 10'b0000000001, 10'b0000000100, 10'b0000001010, 10'b1111110111, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b1111101010, 10'b1111110110, 10'b0000010100, 10'b1111111111, 10'b1111111110, 10'b0000000000, 10'b1111110011, 10'b0000000000, 10'b0000001000, 10'b0000000001, 10'b0000000001, 10'b0000001010, 10'b0000000000, 10'b0000000001, 10'b0000000000, 10'b1111111110, 10'b1111111001, 10'b1111101010, 10'b0000001000, 10'b0000001010, 10'b1111111111, 10'b1111111000, 10'b0000000000, 10'b1111101011, 10'b1111111110, 10'b1111111111, 10'b0000000110, 10'b1111111011, 10'b1111111111, 10'b0000011011, 10'b0000001110, 10'b1111111111, 10'b1111111111, 10'b1111111111, 10'b1111111000, 10'b0000000100, 10'b0000000100, 10'b0000000101, 10'b0000000101, 10'b0000001100, 10'b0000001011, 10'b0000010101, 10'b1111111011, 10'b0000001100, 10'b0000000100, 10'b1111110101, 10'b0000000011, 10'b1111110011, 10'b1111110001, 10'b1111110000}, 
{10'b0000000000, 10'b0000000111, 10'b1111111001, 10'b0000000000, 10'b1111111110, 10'b1111111110, 10'b1111101010, 10'b1111111111, 10'b0000001000, 10'b0000000111, 10'b0000000111, 10'b1111110011, 10'b1111111101, 10'b0000001001, 10'b1111111111, 10'b0000000000, 10'b1111100101, 10'b1111111111, 10'b0000001011, 10'b0000000010, 10'b0000000111, 10'b1111111100, 10'b0000000111, 10'b0000001100, 10'b1111110100, 10'b1111110111, 10'b1111111111, 10'b1111111101, 10'b0000000010, 10'b0000000000, 10'b1111111111, 10'b0000001010, 10'b1111101000, 10'b0000001011, 10'b0000010000, 10'b0000000011, 10'b0000000011, 10'b1111111100, 10'b0000000011, 10'b1111111100, 10'b1111110111, 10'b1111111110, 10'b0000000101, 10'b0000010110, 10'b1111100100, 10'b1111110001, 10'b0000000110, 10'b1111111100, 10'b0000001110, 10'b1111111000, 10'b1111110101, 10'b1111110111, 10'b1111111111, 10'b0000000011, 10'b1111111010, 10'b1111100101, 10'b1111111011, 10'b1111111111, 10'b0000000001, 10'b1111101100, 10'b0000100011, 10'b1111101110, 10'b0000010001, 10'b0000000100}, 
{10'b0000000010, 10'b1111111001, 10'b0000010100, 10'b1111110110, 10'b1111110001, 10'b0000000010, 10'b0000001001, 10'b0000001001, 10'b1111111010, 10'b1111111010, 10'b0000000001, 10'b0000000111, 10'b0000000111, 10'b0000000001, 10'b1111111001, 10'b0000000100, 10'b0000001111, 10'b1111111111, 10'b1111110111, 10'b0000000000, 10'b0000000010, 10'b0000000000, 10'b1111110110, 10'b0000000011, 10'b0000011001, 10'b0000000000, 10'b0000000101, 10'b1111100110, 10'b1111111101, 10'b0000000000, 10'b1111111001, 10'b1111110110, 10'b0000001110, 10'b1111111111, 10'b1111111110, 10'b1111110110, 10'b0000000100, 10'b0000001001, 10'b1111111111, 10'b1111111110, 10'b1111111010, 10'b0000000111, 10'b0000000000, 10'b1111101010, 10'b0000001001, 10'b0000001100, 10'b1111111111, 10'b0000000000, 10'b1111110010, 10'b1111111101, 10'b1111111111, 10'b1111110101, 10'b0000000000, 10'b1111111010, 10'b0000000001, 10'b1111100101, 10'b1111111111, 10'b1111111111, 10'b0000001000, 10'b0000010010, 10'b1111101001, 10'b0000010000, 10'b0000000001, 10'b1111111101}, 
{10'b0000001001, 10'b0000100111, 10'b0000001111, 10'b0000001001, 10'b1111110000, 10'b1111110101, 10'b1110101100, 10'b1111110001, 10'b0000001100, 10'b1111111111, 10'b0000001001, 10'b0000011011, 10'b0000000010, 10'b0000000000, 10'b1111111111, 10'b0000000000, 10'b1111111001, 10'b1111111001, 10'b0000000111, 10'b1111101111, 10'b1111101010, 10'b1111111100, 10'b1111101101, 10'b0000000000, 10'b1110110111, 10'b0000011010, 10'b0000011111, 10'b0000010011, 10'b1111001000, 10'b1111110101, 10'b1111101001, 10'b1111100101, 10'b1110101111, 10'b0000010101, 10'b1111111110, 10'b0000001010, 10'b0000000000, 10'b1111010010, 10'b0000000000, 10'b0000000000, 10'b0000000001, 10'b0000100000, 10'b1111111001, 10'b1111101011, 10'b0000011100, 10'b1111110001, 10'b1111110101, 10'b1111110011, 10'b0000001111, 10'b0000010001, 10'b1111111101, 10'b1111110100, 10'b1111111111, 10'b1111111100, 10'b0000000000, 10'b1111110011, 10'b0000010011, 10'b0000100010, 10'b0000010110, 10'b1111100010, 10'b1110001001, 10'b0000011100, 10'b0000000010, 10'b0000001010}, 
{10'b1111111000, 10'b0000001010, 10'b0000001010, 10'b1111111111, 10'b1111110100, 10'b1111111101, 10'b1111110011, 10'b1111111110, 10'b0000000100, 10'b1111111101, 10'b1111111111, 10'b1111111110, 10'b1111111111, 10'b1111111010, 10'b1111111111, 10'b1111111100, 10'b0000001010, 10'b1111111111, 10'b1111101011, 10'b0000001110, 10'b0000010011, 10'b0000001101, 10'b1111110101, 10'b1111111011, 10'b1111110100, 10'b1111110110, 10'b0000000111, 10'b0000000111, 10'b0000000111, 10'b0000001011, 10'b0000000001, 10'b0000001100, 10'b1111111110, 10'b0000000000, 10'b0000001001, 10'b0000000100, 10'b1111111101, 10'b1111111111, 10'b0000000000, 10'b1111110110, 10'b1111111000, 10'b1111111100, 10'b1111110100, 10'b0000001110, 10'b0000000000, 10'b1111111111, 10'b1111111101, 10'b1111111011, 10'b1111100110, 10'b1111111110, 10'b1111111000, 10'b1111111011, 10'b1111111100, 10'b0000001000, 10'b0000010101, 10'b0000000101, 10'b1111111111, 10'b1111110101, 10'b1111111111, 10'b0000000000, 10'b0000001010, 10'b1111111111, 10'b0000000001, 10'b0000000000}
};

localparam logic signed [9:0] bias [64] = '{
10'b1111111110,  // -0.037350185215473175
10'b0000001000,  // 0.27355897426605225
10'b1111111100,  // -0.12378914654254913
10'b1111111101,  // -0.064457006752491
10'b0000000001,  // 0.05452875792980194
10'b0000000011,  // 0.11671770364046097
10'b0000000100,  // 0.13640816509723663
10'b0000000010,  // 0.07482525706291199
10'b0000000001,  // 0.04674031585454941
10'b1111111001,  // -0.20146161317825317
10'b1111111100,  // -0.09910125285387039
10'b0000000100,  // 0.15104414522647858
10'b1111111100,  // -0.10221704095602036
10'b1111111011,  // -0.1461549550294876
10'b1111111101,  // -0.08641516417264938
10'b0000000101,  // 0.16613510251045227
10'b1111111101,  // -0.0836295336484909
10'b1111111110,  // -0.05756539851427078
10'b1111111110,  // -0.03229188174009323
10'b1111111111,  // -0.028388574719429016
10'b0000000100,  // 0.1260243058204651
10'b1111111110,  // -0.037064336240291595
10'b0000000110,  // 0.19336333870887756
10'b0000000000,  // 0.02124214917421341
10'b0000001111,  // 0.4985624849796295
10'b0000000000,  // 0.0158411655575037
10'b1111111101,  // -0.08296407759189606
10'b0000000011,  // 0.11056788265705109
10'b0000000000,  // 0.01173810102045536
10'b1111111100,  // -0.10843746364116669
10'b0000001000,  // 0.27439257502555847
10'b0000000010,  // 0.09199801832437515
10'b0000001000,  // 0.27419957518577576
10'b0000001000,  // 0.27063727378845215
10'b1111111000,  // -0.24828937649726868
10'b0000000010,  // 0.07818280160427094
10'b1111111111,  // -0.005749030504375696
10'b0000000011,  // 0.10850494354963303
10'b0000000100,  // 0.13591453433036804
10'b1111111100,  // -0.12088628858327866
10'b1111111110,  // -0.05666546896100044
10'b0000000010,  // 0.09311636537313461
10'b0000000001,  // 0.05477767437696457
10'b0000000000,  // 0.029585206881165504
10'b1111110110,  // -0.31209176778793335
10'b1111111101,  // -0.08465463668107986
10'b1111111010,  // -0.16775836050510406
10'b0000000100,  // 0.14762157201766968
10'b1111111000,  // -0.23618532717227936
10'b0000000010,  // 0.06535740196704865
10'b1111111011,  // -0.12853026390075684
10'b1111111011,  // -0.13802281022071838
10'b1111111011,  // -0.15156887471675873
10'b0000000010,  // 0.07979883998632431
10'b0000000101,  // 0.18141601979732513
10'b1111111110,  // -0.054039113223552704
10'b1111111111,  // -0.010052933357656002
10'b0000000010,  // 0.06611225008964539
10'b0000000001,  // 0.05053366720676422
10'b0000000000,  // 0.026860840618610382
10'b0000000001,  // 0.03283466026186943
10'b0000000100,  // 0.15558314323425293
10'b1111110110,  // -0.2863388657569885
10'b1111111101   // -0.08769102394580841
};
endpackage