// Width: 22
// NFRAC: 11
package dense_3_22_11;

localparam logic signed [21:0] weights [32][32] = '{ 
{22'b1111111111111110011011, 22'b1111111111110010000000, 22'b1111111111110011000001, 22'b1111111111111001111001, 22'b0000000000001010111110, 22'b0000000000000001011001, 22'b1111111111111111100101, 22'b1111111111111111111110, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b0000000000000100000010, 22'b1111111111101111001000, 22'b1111111111111110000101, 22'b0000000000011011000110, 22'b1111111111111000010001, 22'b1111111111100010001001, 22'b1111111111111110110101, 22'b0000000000000011100100, 22'b0000000000001101111010, 22'b1111111111110100110110, 22'b1111111111011101111001, 22'b1111111111111110100001, 22'b0000000000000001100100, 22'b1111111111110011000110, 22'b0000000000000000000000, 22'b0000000000100000011001, 22'b1111111111010001011001, 22'b1111111111111000111010, 22'b1111111111110011100100, 22'b1111111111111011001100, 22'b0000000000001101100010, 22'b1111111111111010111001}, 
{22'b0000000000010111111011, 22'b0000000000110111010111, 22'b0000000000001100110111, 22'b1111111111101010111101, 22'b0000000000000111110100, 22'b1111111111110111010000, 22'b1111111111111100100001, 22'b0000000000100010111000, 22'b0000000000000000001100, 22'b1111111111111111111111, 22'b1111111111111110111110, 22'b1111111111101101001011, 22'b1111111111111001100011, 22'b0000000000010001010010, 22'b1111111110111100100111, 22'b1111111111110000111010, 22'b1111111111111111111111, 22'b1111111111111111101111, 22'b1111111111111110010100, 22'b1111111111111010101111, 22'b1111111111110111101110, 22'b1111111111110111001100, 22'b0000000000000000100011, 22'b1111111111111111111100, 22'b1111111111111111110010, 22'b1111111111011101101100, 22'b0000000000000000011000, 22'b0000000000001111000100, 22'b1111111111111101111110, 22'b1111111111101001111011, 22'b0000000000000000000101, 22'b0000000000000001001101}, 
{22'b1111111111100000011110, 22'b0000000000000101111001, 22'b0000000000000000010101, 22'b0000000000001010010100, 22'b1111111111101011110101, 22'b0000000000000000000001, 22'b0000000000000000000011, 22'b1111111111100101001001, 22'b0000000000010001001001, 22'b1111111111110111100111, 22'b1111111111110111101100, 22'b1111111111010000011010, 22'b1111111111110110000011, 22'b0000000000010000010110, 22'b0000000000001000011100, 22'b1111111111111111111100, 22'b1111111111111100010101, 22'b1111111111111111001111, 22'b1111111111100101111011, 22'b0000000000000000000110, 22'b0000000000000011111111, 22'b0000000000000010001101, 22'b0000000000000110101100, 22'b0000000000011100001010, 22'b0000000000000001001101, 22'b1111111111100110110001, 22'b0000000000011000100011, 22'b0000000000000000000001, 22'b0000000000000101010011, 22'b1111111111111111010010, 22'b0000000000000000000001, 22'b0000000001001000100110}, 
{22'b0000000000011010110011, 22'b1111111111111111111111, 22'b1111111111111001110001, 22'b0000000000101001111000, 22'b0000000000100111010011, 22'b0000000000000000000000, 22'b0000000000000010010110, 22'b0000000000011010000010, 22'b1111111111110011010101, 22'b1111111111111111111111, 22'b1111111111100101101001, 22'b0000000000000011110101, 22'b0000000000001000100001, 22'b1111111111101000000101, 22'b0000000000000010111111, 22'b1111111111111010111000, 22'b1111111111111111111111, 22'b1111111111110100010110, 22'b0000000000000001001110, 22'b0000000000000001110001, 22'b0000000000000000100000, 22'b1111111111111101101010, 22'b0000000000100110001100, 22'b0000000000010101111100, 22'b0000000000010101000101, 22'b0000000000001111111000, 22'b0000000000010101110111, 22'b0000000000000000000000, 22'b1111111111111100001110, 22'b0000000000011100111111, 22'b0000000000001111111110, 22'b1111111111111010011000}, 
{22'b0000000000100000000001, 22'b1111111111111101000000, 22'b1111111111101001110100, 22'b1111111111001111111001, 22'b0000000000011110100011, 22'b0000000000000000000000, 22'b1111111111100101101111, 22'b1111111111101101111010, 22'b1111111111111101000001, 22'b1111111111001100001101, 22'b1111111110111001010010, 22'b0000000000011110010000, 22'b0000000000101010110011, 22'b0000000000100001011111, 22'b1111111111011011001100, 22'b1111111111001110011001, 22'b0000000000000000000000, 22'b1111111111110110111100, 22'b0000000000001100110110, 22'b0000000000001000111000, 22'b1111111111110011111100, 22'b1111111111111111100101, 22'b0000000000101110001011, 22'b1111111110101000000001, 22'b0000000000000101101000, 22'b1111111111010101110110, 22'b0000000000000100001100, 22'b1111111111110000000111, 22'b1111111111101100111001, 22'b1111111111111111111110, 22'b0000000000000100011110, 22'b0000000000100101001001}, 
{22'b0000000000000010110000, 22'b1111111111111101010110, 22'b1111111111101100010110, 22'b1111111111101111010101, 22'b0000000000010111110010, 22'b0000000000000000000000, 22'b1111111111101110000110, 22'b1111111111110111010010, 22'b1111111111100100100110, 22'b1111111111111011111001, 22'b1111111111111111111110, 22'b0000000000001010010000, 22'b0000000000000000000000, 22'b0000000000010110111001, 22'b1111111111011111101000, 22'b1111111111110111110101, 22'b0000000000000101101100, 22'b1111111111101101001111, 22'b1111111111110011010110, 22'b1111111111111111111111, 22'b0000000000000000110001, 22'b0000000000010011001011, 22'b0000000000011101111000, 22'b1111111111111111010100, 22'b1111111111111111111110, 22'b0000000000011001101001, 22'b1111111111011100110101, 22'b1111111111111111111111, 22'b1111111111110000110111, 22'b1111111111111101101001, 22'b1111111111111111110011, 22'b0000000000000000011010}, 
{22'b0000000000000100001010, 22'b1111111111101010101110, 22'b0000000000000110111011, 22'b1111111111111101100010, 22'b1111111111111111100001, 22'b0000000000001001101100, 22'b1111111111111001001101, 22'b1111111111010100101010, 22'b1111111111111111111111, 22'b1111111111110010101010, 22'b1111111111100010110001, 22'b0000000000011110001110, 22'b0000000000000000011101, 22'b0000000000101011110011, 22'b0000000000110101000010, 22'b0000000000000000001010, 22'b1111111111111111111111, 22'b1111111111101011110100, 22'b1111111111111100000010, 22'b0000000000010001011111, 22'b1111111111001111111111, 22'b0000000000001001111110, 22'b0000000000010100111000, 22'b0000000000000001001101, 22'b0000000000001001100110, 22'b0000000001001111100100, 22'b1111111111100110110001, 22'b1111111111111010001100, 22'b1111111111110011110110, 22'b0000000000011111001011, 22'b1111111111111100110110, 22'b1111111111110101001010}, 
{22'b1111111111011001110101, 22'b0000000000000001100001, 22'b1111111111010111101110, 22'b0000000000011011110110, 22'b0000000001000001110010, 22'b0000000000000111011011, 22'b0000000000000000001111, 22'b0000000000000011000001, 22'b1111111111111111111111, 22'b0000000000001000001100, 22'b0000000001010011010001, 22'b1111111111111111111110, 22'b0000000000011000011001, 22'b0000000000100111110111, 22'b0000000000110001001100, 22'b0000000001000011001101, 22'b0000000000000000000000, 22'b1111111111100001011001, 22'b0000000000010101100001, 22'b1111111111111111101001, 22'b1111111111010111001011, 22'b1111111111110001011110, 22'b0000000000000000110111, 22'b1111111111111010101100, 22'b1111111111011111111010, 22'b0000000001111000000010, 22'b1111111111110001111100, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b0000000000111000100000, 22'b0000000000000101101011, 22'b0000000000011001000100}, 
{22'b0000000000011011000001, 22'b1111111111111110110000, 22'b0000000000000000000001, 22'b1111111111111101001110, 22'b0000000000000101001110, 22'b1111111111111101100100, 22'b1111111111111111111110, 22'b0000000000001010000010, 22'b0000000000001101100001, 22'b1111111111101110011101, 22'b0000000000001000111101, 22'b0000000000001011111111, 22'b0000000000000000110000, 22'b0000000000010101010011, 22'b1111111111110001100110, 22'b1111111111001100111111, 22'b0000000000000000000000, 22'b1111111111111111000110, 22'b1111111111111110010010, 22'b1111111111100000000101, 22'b1111111111111111111011, 22'b0000000000000000000000, 22'b1111111111110011000001, 22'b1111111111111111000110, 22'b1111111111111001111010, 22'b0000000000001001111110, 22'b0000000000010111111010, 22'b1111111111111000010110, 22'b1111111111111100110110, 22'b1111111111111101011011, 22'b0000000000000001101110, 22'b1111111111100110111000}, 
{22'b1111111111110100101000, 22'b0000000000011000100110, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b0000000000110010101101, 22'b0000000000010100100111, 22'b1111111111111111111111, 22'b1111111111011100011110, 22'b0000000000000111100010, 22'b1111111111010011010110, 22'b1111111110100110001100, 22'b1111111111111111111111, 22'b0000000000000000000001, 22'b0000000000011011011101, 22'b0000000000000111000110, 22'b0000000000000000000000, 22'b1111111111101010111110, 22'b0000000000000000000001, 22'b0000000000000000011011, 22'b0000000000000011111000, 22'b0000000000001111100110, 22'b1111111111111110010111, 22'b1111111111101000111100, 22'b0000000000000000100001, 22'b1111111111111111010001, 22'b0000000001000101001101, 22'b0000000000010100111001, 22'b1111111111111111111110, 22'b1111111111111011011101, 22'b0000000000101010110001, 22'b1111111111111101011100, 22'b1111111111111010011001}, 
{22'b1111111111011110100001, 22'b0000000000001011001101, 22'b1111111111111101110001, 22'b1111111111111111111111, 22'b1111111111110000001111, 22'b1111111111100111110101, 22'b0000000000000011000100, 22'b0000000000001001001110, 22'b1111111111111111111111, 22'b1111111111110101000010, 22'b1111111111011011010110, 22'b0000000000001100110110, 22'b0000000000010011011101, 22'b0000000000000000000000, 22'b0000000000110101101100, 22'b1111111111011100000011, 22'b0000000000000110101001, 22'b1111111111100110111110, 22'b0000000000010010000011, 22'b1111111111111111111111, 22'b1111111111111101100010, 22'b0000000000000100011111, 22'b0000000000000111110110, 22'b0000000000000000000000, 22'b1111111111100000011001, 22'b0000000000000001111111, 22'b1111111111011100001111, 22'b1111111111111101011101, 22'b1111111111111111111111, 22'b0000000000101011001111, 22'b1111111111110011110101, 22'b0000000000000000000001}, 
{22'b1111111111111111111111, 22'b0000000000000111010110, 22'b0000000000000000000001, 22'b0000000000011001000010, 22'b1111111111111000100000, 22'b1111111111111101001111, 22'b0000000000000011101111, 22'b1111111111111111101000, 22'b1111111111111101000010, 22'b0000000000101001000000, 22'b0000000000101100101111, 22'b0000000000000000000010, 22'b1111111111101010101101, 22'b1111111111010011000011, 22'b1111111111111100110000, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b1111111111111011111011, 22'b1111111111100001100000, 22'b0000000000011000011110, 22'b0000000000000000001000, 22'b0000000000010111101111, 22'b1111111111111111111111, 22'b0000000000100011111111, 22'b0000000000000111111010, 22'b0000000000010011100110, 22'b0000000000011101001001, 22'b1111111111111100101100, 22'b1111111111100110111100, 22'b1111111111100011110011, 22'b1111111111111111101011, 22'b1111111111010101001100}, 
{22'b1111111111110001100000, 22'b1111111111111111111111, 22'b0000000000000111101000, 22'b1111111111100101001100, 22'b0000000000000101100000, 22'b1111111111111111111111, 22'b1111111111110010000110, 22'b1111111111111111011000, 22'b1111111111110111111110, 22'b0000000000000010011000, 22'b0000000000000100111111, 22'b1111111111111011011011, 22'b0000000000000001000011, 22'b0000000000001100000000, 22'b1111111111010111111111, 22'b1111111111110000010101, 22'b0000000000001110100110, 22'b1111111111110100101011, 22'b0000000000000000000000, 22'b1111111111111110011001, 22'b0000000000001100010110, 22'b0000000000000000100000, 22'b1111111111111110000000, 22'b0000000000000010101110, 22'b0000000000010001001111, 22'b1111111111111001010110, 22'b0000000000000000000000, 22'b1111111111100011000101, 22'b1111111111110011011110, 22'b1111111111111111100011, 22'b0000000000001011000110, 22'b0000000000000000000001}, 
{22'b1111111111011110101111, 22'b0000000000011010111001, 22'b1111111111111111111111, 22'b1111111111111111100100, 22'b1111111111111111011000, 22'b0000000000001011001110, 22'b1111111111111111111111, 22'b0000000000110001011010, 22'b1111111111111111000011, 22'b1111111111111111111111, 22'b0000000000001101001011, 22'b0000000000000010100111, 22'b0000000000000000011010, 22'b0000000000000000000000, 22'b0000000000000111110010, 22'b0000000000010101001000, 22'b0000000000001011011001, 22'b0000000000001010101010, 22'b1111111111111111011101, 22'b0000000000010011101010, 22'b0000000000000110011100, 22'b0000000000000010100101, 22'b1111111111111111011100, 22'b0000000000010000010000, 22'b1111111111111001101000, 22'b1111111111101010010011, 22'b1111111111111010000101, 22'b1111111111111111111111, 22'b0000000000000110100000, 22'b0000000000000001111001, 22'b0000000000001100100000, 22'b0000000000011110101010}, 
{22'b1111111111111110110011, 22'b1111111111100111000101, 22'b0000000000000011010011, 22'b1111111111111111111100, 22'b0000000000111010101000, 22'b1111111111110010101110, 22'b1111111111011011011010, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b1111111111111110010110, 22'b0000000000000011000110, 22'b0000000000011011111100, 22'b0000000000010100100110, 22'b0000000000000000101011, 22'b0000000000000010001000, 22'b1111111111110100110100, 22'b0000000000000010001000, 22'b1111111111111101100100, 22'b0000000000000000000000, 22'b0000000000000100110100, 22'b1111111111111101100110, 22'b0000000000000001001110, 22'b0000000000010001000010, 22'b0000000000000010010111, 22'b1111111111111111001110, 22'b1111111111100101100101, 22'b0000000000001101000000, 22'b1111111111111111111111, 22'b1111111111111111111110, 22'b1111111111111001001100, 22'b1111111111111110101000, 22'b1111111111111011111111}, 
{22'b0000000000000000011101, 22'b1111111111111011111100, 22'b1111111111110111111011, 22'b1111111111110010000000, 22'b1111111111011101000001, 22'b0000000000100111000000, 22'b0000000000000000000000, 22'b0000000000001010110011, 22'b0000000000010010010111, 22'b0000000000000000110100, 22'b1111111111111101110101, 22'b0000000000011110011100, 22'b0000000000001110010100, 22'b1111111111101000100110, 22'b1111111111110101100111, 22'b1111111111111101010111, 22'b1111111111100110100000, 22'b1111111111111110111000, 22'b0000000000000000000000, 22'b1111111111111111101101, 22'b0000000000001001111110, 22'b1111111111110111001111, 22'b0000000000000000000000, 22'b0000000000000100111011, 22'b1111111111111111111111, 22'b1111111111101010001000, 22'b0000000000001010000001, 22'b0000000000000000000001, 22'b0000000000000010110110, 22'b0000000000000000101100, 22'b1111111111101011110001, 22'b0000000000000001010101}, 
{22'b1111111111110011011100, 22'b1111111111110101111011, 22'b0000000000000100111001, 22'b1111111111111000000011, 22'b1111111111111010010000, 22'b0000000000000111011011, 22'b1111111111111111101011, 22'b0000000000000010001111, 22'b0000000000001000011000, 22'b1111111111111111111110, 22'b0000000000000111111010, 22'b1111111111110111110110, 22'b1111111111111111011000, 22'b1111111111111111111111, 22'b0000000000000110100111, 22'b1111111111111111111111, 22'b0000000000011111010000, 22'b1111111111111110111000, 22'b0000000000001111111000, 22'b1111111111110101001000, 22'b0000000000001010001000, 22'b0000000000000100000001, 22'b0000000000000101011001, 22'b0000000000000010010100, 22'b1111111111111010110010, 22'b1111111111101110001010, 22'b1111111111101111011010, 22'b0000000000000110111010, 22'b1111111111111010101001, 22'b0000000000000000000010, 22'b1111111111111110001111, 22'b0000000000001110110110}, 
{22'b1111111111111111111111, 22'b1111111111100110000101, 22'b1111111111100110100111, 22'b1111111111111111111111, 22'b0000000000101000011001, 22'b1111111111111010001100, 22'b0000000000000000000000, 22'b0000000000011110111011, 22'b1111111111110110100011, 22'b0000000000000000000000, 22'b1111111111100101010001, 22'b1111111111100000101000, 22'b0000000000011100101100, 22'b0000000000001001101011, 22'b1111111111111000001111, 22'b1111111111101110011110, 22'b0000000000001011000010, 22'b0000000000000000000001, 22'b1111111111110000110010, 22'b0000000000000001101100, 22'b0000000000000100011100, 22'b1111111111111010010101, 22'b0000000000010010001011, 22'b1111111111000001010011, 22'b0000000000000010100111, 22'b0000000000001111010011, 22'b1111111111111101010111, 22'b0000000000000000111101, 22'b1111111111110001000100, 22'b1111111111111111111111, 22'b1111111111110011001000, 22'b1111111111111110011101}, 
{22'b0000000000001101100110, 22'b0000000000010110000101, 22'b0000000000100011001111, 22'b1111111111110010111010, 22'b0000000000011010101000, 22'b0000000000010011100110, 22'b0000000000000000000010, 22'b0000000000011101001001, 22'b0000000000010110110110, 22'b1111111111111001001010, 22'b0000000000101100111001, 22'b1111111111101001101001, 22'b0000000000100111110001, 22'b0000000000011100100100, 22'b1111111110111011010101, 22'b1111111111111111111100, 22'b0000000000000000000000, 22'b0000000000000000010111, 22'b0000000000010000101000, 22'b1111111111011111110010, 22'b0000000000001110001011, 22'b1111111111110010011011, 22'b1111111111100000100111, 22'b1111111111110101111101, 22'b0000000000010101000101, 22'b1111111111010101110001, 22'b1111111111101010111001, 22'b1111111111111101010111, 22'b1111111111111111111111, 22'b1111111111011011111000, 22'b0000000000011001010011, 22'b0000000000000000000001}, 
{22'b1111111111111100110110, 22'b0000000000000000000010, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b1111111111101001100001, 22'b0000000000000000100101, 22'b0000000000000000100001, 22'b1111111111111111000010, 22'b1111111111111110011100, 22'b1111111111111101000011, 22'b0000000000001000111001, 22'b1111111111111111111100, 22'b0000000000000101010011, 22'b1111111111101010000110, 22'b0000000000000110110101, 22'b1111111111111111111101, 22'b0000000000001001000000, 22'b0000000000011100101001, 22'b1111111111101001011011, 22'b0000000000000011010100, 22'b1111111111111001101010, 22'b0000000000001000001110, 22'b0000000000001100001010, 22'b1111111111111010100010, 22'b1111111111101111111011, 22'b0000000000000001010100, 22'b0000000000110101000100, 22'b1111111111111110011100, 22'b1111111111111111000001, 22'b0000000000010100110000, 22'b0000000000000000000000, 22'b0000000000110111001010}, 
{22'b1111111111011110100111, 22'b0000000000000010010100, 22'b1111111111110010001001, 22'b0000000000011000100000, 22'b0000000000000111000001, 22'b1111111111111101111110, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b1111111111101100100110, 22'b1111111111111101111000, 22'b0000000000000000000000, 22'b1111111111011100011101, 22'b0000000000000000110011, 22'b1111111111111101011101, 22'b1111111111111111110101, 22'b1111111111111111111111, 22'b1111111111111000100010, 22'b0000000000000000010110, 22'b0000000000000000001100, 22'b0000000000001010001001, 22'b0000000000000001000111, 22'b0000000000000000000000, 22'b0000000000000000000000, 22'b1111111111111111011110, 22'b0000000000000000000001, 22'b0000000000000001001011, 22'b0000000000100101001101, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b1111111111111101011001, 22'b0000000000001011001101, 22'b1111111111111110010111}, 
{22'b1111111111111111111001, 22'b1111111111110110010100, 22'b0000000000001101000100, 22'b0000000000000010100011, 22'b1111111111101000001101, 22'b0000000000000000000010, 22'b0000000000010010010011, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b1111111111111001101100, 22'b0000000000000111010110, 22'b0000000000000001001101, 22'b0000000000010100101101, 22'b1111111111011100111010, 22'b1111111111111001111100, 22'b1111111111111110111001, 22'b0000000000001101110101, 22'b1111111111100111011010, 22'b0000000000000001010111, 22'b1111111111001111101101, 22'b1111111111111110110010, 22'b1111111111111000011000, 22'b1111111111111101011010, 22'b0000000000010010111011, 22'b1111111111111011001110, 22'b1111111111101110000000, 22'b0000000000000101110010, 22'b0000000000000000000001, 22'b0000000000011001010101, 22'b0000000000100001011111, 22'b1111111111101011000000, 22'b1111111111100011010000}, 
{22'b0000000000000100010100, 22'b0000000000000001101000, 22'b1111111111100101011111, 22'b1111111111111100010111, 22'b1111111111111111111111, 22'b0000000000000000001000, 22'b0000000000000110110011, 22'b0000000000011010010100, 22'b0000000000000000000000, 22'b0000000000000001010011, 22'b0000000000000100011110, 22'b1111111111011101011110, 22'b1111111111111011101111, 22'b1111111111011001010111, 22'b0000000000011110110001, 22'b0000000000000000000001, 22'b1111111111111111111100, 22'b1111111111010110111111, 22'b1111111111111111111110, 22'b1111111111111011001111, 22'b1111111111111110101010, 22'b0000000000000000000000, 22'b0000000000000011111111, 22'b1111111111110110011000, 22'b0000000000000011011001, 22'b0000000000011010010011, 22'b0000000000011011010010, 22'b0000000000011000111111, 22'b0000000000010011101101, 22'b0000000000000000000000, 22'b0000000000000111010011, 22'b0000000000110010001001}, 
{22'b1111111111111110011000, 22'b1111111111110000110001, 22'b0000000000011000111010, 22'b1111111111111001011010, 22'b0000000000000100011101, 22'b0000000000001010101111, 22'b1111111111111111111111, 22'b1111111111101101101000, 22'b1111111111111010100011, 22'b1111111111011001100011, 22'b0000000000011100101000, 22'b0000000000000000001111, 22'b0000000000011010110100, 22'b0000000000101010111000, 22'b1111111111111000100011, 22'b1111111111001000010001, 22'b1111111111111001010110, 22'b0000000000011110000100, 22'b1111111111101101111001, 22'b1111111111110010101001, 22'b0000000000000011110011, 22'b0000000000000000000100, 22'b1111111111011101000111, 22'b1111111111110011110000, 22'b1111111111111101011111, 22'b1111111111111000001101, 22'b0000000000000111001011, 22'b0000000000101101000001, 22'b0000000000001111101101, 22'b1111111111111111111111, 22'b0000000000000101001010, 22'b0000000000000001110001}, 
{22'b0000000000000010101101, 22'b0000000000011101000010, 22'b0000000000000000000000, 22'b0000000000010010111010, 22'b0000000000110101001100, 22'b1111111111110101000100, 22'b1111111111111111111111, 22'b1111111111111101001010, 22'b0000000000010010110000, 22'b1111111111110011101111, 22'b1111111111111111111010, 22'b0000000000010101010101, 22'b0000000000000000100010, 22'b0000000000000001110000, 22'b1111111110011110010001, 22'b1111111111111010111010, 22'b0000000000000000000000, 22'b0000000000001100110110, 22'b1111111111111111110010, 22'b0000000000010011000111, 22'b1111111111111111111111, 22'b1111111111110100111100, 22'b1111111111011100000010, 22'b0000000000001000010111, 22'b0000000000010010010011, 22'b1111111110111001000000, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b0000000000100010110100, 22'b1111111111001100101101, 22'b0000000000000000000111, 22'b1111111111111111100111}, 
{22'b0000000000000000100110, 22'b1111111111101010010000, 22'b0000000000000011011101, 22'b1111111111111111000010, 22'b0000000000000011010101, 22'b0000000000100001110111, 22'b1111111111010001100111, 22'b0000000000000010001100, 22'b0000000000011011000110, 22'b1111111111101010011010, 22'b1111111111111110100000, 22'b0000000000000011001000, 22'b1111111111111111011011, 22'b0000000000001011011100, 22'b0000000000000110110111, 22'b1111111111111110111011, 22'b0000000000000100010010, 22'b0000000000000000000001, 22'b0000000000000001011000, 22'b0000000000011000010011, 22'b1111111111111110001101, 22'b1111111111100001000000, 22'b1111111111011001010010, 22'b1111111111110011100110, 22'b1111111111011010001100, 22'b0000000000001101010100, 22'b0000000000100111111000, 22'b0000000000010111100110, 22'b1111111111111111010101, 22'b1111111111101000001001, 22'b1111111111101100000111, 22'b0000000000000011110100}, 
{22'b0000000000000011010100, 22'b1111111111100001011011, 22'b1111111111111110111010, 22'b0000000000001001101000, 22'b1111111111100001011000, 22'b0000000000001010110111, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b0000000000000000000000, 22'b0000000000010000111010, 22'b1111111111111110111001, 22'b0000000000000000100111, 22'b0000000000000000000001, 22'b0000000000001000001001, 22'b1111111111111110111010, 22'b0000000000000000001011, 22'b1111111111111111111101, 22'b1111111111101011011000, 22'b1111111111011111101000, 22'b1111111111111111111101, 22'b1111111111011101110101, 22'b1111111111101100101110, 22'b1111111111101000001101, 22'b0000000000111000111111, 22'b0000000000000001001000, 22'b1111111111111101000011, 22'b0000000000010100010011, 22'b0000000000111001011100, 22'b0000000000011001010001, 22'b1111111110111100001000, 22'b1111111111110100001000}, 
{22'b0000000000011000000011, 22'b1111111111111111111110, 22'b0000000000010000000100, 22'b1111111111111110101110, 22'b0000000000011110111101, 22'b1111111111110110110111, 22'b0000000000000100100010, 22'b0000000000011010110001, 22'b0000000000010001001000, 22'b1111111111011110100101, 22'b1111111111111100000011, 22'b0000000000000111110111, 22'b0000000000000100011010, 22'b1111111111111111000100, 22'b0000000000000101011011, 22'b0000000000000000000001, 22'b0000000000010111001100, 22'b0000000000000010001111, 22'b0000000000010111111100, 22'b1111111111111011110011, 22'b1111111111110111110110, 22'b1111111111111011001101, 22'b1111111111111111111111, 22'b0000000000010011010100, 22'b1111111111110011000011, 22'b1111111111111111100110, 22'b0000000000000000000000, 22'b0000000000000000000001, 22'b0000000000000000000000, 22'b0000000000010010101100, 22'b1111111111101011011110, 22'b1111111111111110100000}, 
{22'b1111111111111111111101, 22'b1111111111111110000001, 22'b1111111111100010001111, 22'b0000000000010010001101, 22'b0000000000001110010010, 22'b1111111111111000111111, 22'b1111111111111111111111, 22'b1111111111110001011110, 22'b0000000000000000011011, 22'b1111111111111111111110, 22'b1111111111101100101101, 22'b1111111111110000001111, 22'b0000000000011110101010, 22'b0000000000000000000000, 22'b1111111111110111110100, 22'b1111111111111111111111, 22'b0000000000001101101100, 22'b1111111111111111111111, 22'b1111111111111111111111, 22'b1111111111110010001011, 22'b0000000000010100001111, 22'b0000000000000000000000, 22'b0000000000001001111111, 22'b1111111111111110001010, 22'b0000000000001010000011, 22'b0000000000000000001001, 22'b0000000000000000000000, 22'b0000000000001111011010, 22'b1111111111110011101101, 22'b1111111111111101000011, 22'b0000000000001010010001, 22'b1111111111111001001110}, 
{22'b1111111111111110111011, 22'b1111111111101100010000, 22'b0000000000100110000010, 22'b1111111111111011110101, 22'b0000000000001100100100, 22'b1111111111101101101100, 22'b0000000000000000000000, 22'b0000000000000010001100, 22'b1111111111100001010101, 22'b1111111111111111001011, 22'b1111111111111000000101, 22'b0000000000000011101110, 22'b1111111111101011000000, 22'b0000000000001000110100, 22'b0000000000001100111100, 22'b0000000000000111000000, 22'b0000000000000101011111, 22'b1111111111111101100100, 22'b1111111111010010101011, 22'b1111111111111111001000, 22'b1111111111111100010110, 22'b0000000000001000111100, 22'b1111111111111000111001, 22'b1111111111111111111111, 22'b0000000000001100101001, 22'b1111111111111101000101, 22'b1111111111111111000100, 22'b0000000000011000111001, 22'b1111111111100110100001, 22'b1111111111101101000111, 22'b0000000000010110011100, 22'b0000000000000010010011}, 
{22'b0000000000011011100101, 22'b0000000000001100111000, 22'b0000000000000000000011, 22'b1111111111110101110100, 22'b1111111111111010111110, 22'b1111111111111111111100, 22'b0000000000000000000000, 22'b1111111111111011100100, 22'b1111111111111000000011, 22'b1111111111111000011010, 22'b0000000000000000000001, 22'b0000000000001010001000, 22'b0000000000000000011010, 22'b0000000000000011011000, 22'b1111111111111101001001, 22'b0000000000000000010111, 22'b1111111111110110001011, 22'b0000000000000000000010, 22'b1111111111111110110111, 22'b1111111111111111111101, 22'b0000000000000000001001, 22'b0000000000000011110011, 22'b0000000000000110001110, 22'b0000000000000000000000, 22'b0000000000000000000001, 22'b1111111111011000111011, 22'b1111111111110011001111, 22'b0000000000000000011011, 22'b0000000000000001010011, 22'b0000000000000000000101, 22'b1111111111110100101010, 22'b0000000000000001010111}, 
{22'b0000000000001100000000, 22'b1111111110111101001001, 22'b1111111111111111111111, 22'b1111111111111011001011, 22'b1111111111110001000110, 22'b1111111111111111011000, 22'b0000000000000000000000, 22'b0000000000100011000011, 22'b1111111111111101001100, 22'b1111111111111110100110, 22'b0000000000000101010001, 22'b1111111111010101101101, 22'b0000000000000001100010, 22'b1111111111100011111100, 22'b0000000000101110001111, 22'b1111111111111100101001, 22'b1111111111110001100000, 22'b1111111111011100111111, 22'b1111111111111111010100, 22'b1111111111010010101100, 22'b1111111111001100001011, 22'b1111111111111111111110, 22'b0000000000000000000001, 22'b0000000000000000000000, 22'b0000000000001111100111, 22'b1111111111111111000110, 22'b1111111111101100111010, 22'b1111111111111011010110, 22'b1111111111111110100000, 22'b0000000000000000000000, 22'b1111111111111101111110, 22'b1111111111010011001101}
};

localparam logic signed [21:0] bias [32] = '{
22'b0000000000010000111001,  // 0.5280959606170654
22'b0000000000011010111011,  // 0.8414360880851746
22'b0000000000001100101110,  // 0.397830605506897
22'b0000000000001101001000,  // 0.4105983078479767
22'b1111111110001010111100,  // -3.657735586166382
22'b1111111111100011010001,  // -0.8977976441383362
22'b0000000000110110100100,  // 1.7051936388015747
22'b1111111111010111001001,  // -1.2765135765075684
22'b1111111111101101010100,  // -0.5837795734405518
22'b0000000001010110011000,  // 2.699671983718872
22'b0000000000000110111100,  // 0.2170683741569519
22'b0000000000011100001101,  // 0.8814588785171509
22'b1111111110101011101100,  // -2.634300947189331
22'b1111111111000011111011,  // -1.877297282218933
22'b0000000000110101001100,  // 1.6625694036483765
22'b0000000001010111110111,  // 2.7459704875946045
22'b1111111111110000101100,  // -0.47838035225868225
22'b0000000000110110010110,  // 1.6984987258911133
22'b0000000000011011010110,  // 0.8548859357833862
22'b0000000000100000001001,  // 1.0045719146728516
22'b0000000000101101011011,  // 1.4197649955749512
22'b0000000000011010101000,  // 0.832463800907135
22'b0000000000010001011000,  // 0.5434179306030273
22'b0000000000011101101011,  // 0.9277304410934448
22'b1111111111110101000010,  // -0.3426123857498169
22'b1111111111101110000111,  // -0.5587119460105896
22'b1111111111101100001000,  // -0.6208624839782715
22'b1111111111010111000010,  // -1.2802538871765137
22'b0000000000000001111001,  // 0.05940237268805504
22'b1111111111100101101101,  // -0.8213341236114502
22'b0000000000011100000110,  // 0.8783953189849854
22'b1111111111100001100111   // -0.949700653553009
};
endpackage