// Width: 14
// NFRAC: 7
package dense_2_14_7;

localparam logic signed [13:0] weights [64][32] = '{ 
{14'b00000000100010, 14'b00000000000001, 14'b11111111100111, 14'b11111111111101, 14'b00000000100001, 14'b00000000000000, 14'b11111111101101, 14'b11111111111111, 14'b11111111011100, 14'b00000000001010, 14'b00000000000000, 14'b11111111111111, 14'b11111111111111, 14'b11111111100110, 14'b11111111111001, 14'b11111111011110, 14'b00000000000000, 14'b11111111111110, 14'b11111111100111, 14'b11111111101011, 14'b00000000000000, 14'b00000000000000, 14'b11111111111110, 14'b11111111111111, 14'b00000000000000, 14'b00000000001100, 14'b00000000110001, 14'b00000000010110, 14'b11111111111111, 14'b00000000000110, 14'b11111111001011, 14'b00000000000000}, 
{14'b11111111110011, 14'b11111111101100, 14'b11111111101110, 14'b11111111111000, 14'b11111111111111, 14'b00000000000101, 14'b11111111100011, 14'b00000000000000, 14'b00000000000000, 14'b11111111110111, 14'b00000000010011, 14'b11111111111010, 14'b11111111111000, 14'b11111111100100, 14'b00000000000000, 14'b11111111111001, 14'b00000000000001, 14'b11111111100111, 14'b00000000010101, 14'b00000000011101, 14'b11111111111011, 14'b11111111111111, 14'b11111111111111, 14'b00000000000011, 14'b11111111110110, 14'b00000000100011, 14'b00000000011111, 14'b00000000000001, 14'b00000000000011, 14'b11111111000001, 14'b00000000000000, 14'b00000000000000}, 
{14'b00000000001001, 14'b11111111110001, 14'b11111111101111, 14'b11111111111010, 14'b11111111110110, 14'b11111111110101, 14'b11111111101000, 14'b00000000000000, 14'b11111111101110, 14'b00000000000001, 14'b00000000000000, 14'b11111111110101, 14'b00000000001011, 14'b11111111110111, 14'b11111111111111, 14'b11111111111011, 14'b00000000000000, 14'b00000000001100, 14'b00000000000111, 14'b00000000011101, 14'b00000000000101, 14'b11111111110101, 14'b00000000000000, 14'b00000000000100, 14'b11111111111101, 14'b00000000011010, 14'b00000000010011, 14'b00000000001100, 14'b11111111111111, 14'b11111111101100, 14'b11111111111110, 14'b00000000001100}, 
{14'b00000000010001, 14'b00000000000010, 14'b00000000000110, 14'b11111111111110, 14'b11111110111110, 14'b00000000000000, 14'b00000000000000, 14'b00000000011100, 14'b00000000011111, 14'b11111111111110, 14'b11111111111111, 14'b00000000000000, 14'b00000000000000, 14'b00000000000000, 14'b11111111111101, 14'b00000000011011, 14'b00000000000000, 14'b11111111111100, 14'b11111111111111, 14'b11111111101001, 14'b11111111111000, 14'b00000000000110, 14'b11111111110111, 14'b11111111111111, 14'b00000000000000, 14'b11111111111001, 14'b00000000001001, 14'b11111111111111, 14'b11111111111111, 14'b11111111111111, 14'b11111111100100, 14'b00000000100111}, 
{14'b11111110101000, 14'b11111111111100, 14'b11111111111111, 14'b00000000000000, 14'b11111111111100, 14'b00000000000000, 14'b11111111111001, 14'b11111111101100, 14'b00000000000110, 14'b11111111111101, 14'b11111111111110, 14'b11111111111111, 14'b11111111111111, 14'b00000000011010, 14'b00000000000000, 14'b00000000101010, 14'b11111111111111, 14'b00000000011011, 14'b11111111001100, 14'b00000000000000, 14'b11111111110001, 14'b00000000010101, 14'b00000000100001, 14'b00000000000000, 14'b00000000000101, 14'b00000000010100, 14'b00000000011110, 14'b00000000000010, 14'b11111111111111, 14'b11111111111111, 14'b11111111111110, 14'b00000000011100}, 
{14'b00000000000111, 14'b11111111111111, 14'b00000000010011, 14'b11111110101100, 14'b11111101001111, 14'b11111111010011, 14'b00000000101101, 14'b11111110110000, 14'b11111111111111, 14'b11111110101001, 14'b11111110111111, 14'b11111111010100, 14'b00000000101101, 14'b11111111111111, 14'b11111111111110, 14'b00000000000000, 14'b11111111111111, 14'b11111111111111, 14'b11111111101111, 14'b11111111111111, 14'b11111111000001, 14'b00000000000000, 14'b00000000010111, 14'b11111111111111, 14'b00000000000010, 14'b00000000100010, 14'b00000000000110, 14'b11111111111111, 14'b11111111111111, 14'b00000000011010, 14'b11111111111011, 14'b00000000011001}, 
{14'b11111111111011, 14'b11111111101011, 14'b11111111100001, 14'b11111111111001, 14'b11111111011011, 14'b00000000001000, 14'b11111111101000, 14'b11111111101101, 14'b11111111001010, 14'b00000000000110, 14'b11111111111111, 14'b11111111101011, 14'b00000000001111, 14'b11111111111110, 14'b11111111111010, 14'b11111110111001, 14'b11111111111111, 14'b00000000001010, 14'b00000000011000, 14'b11111111101011, 14'b11111111101100, 14'b11111111110111, 14'b11111111111111, 14'b00000000000011, 14'b11111111111010, 14'b11111110101101, 14'b11111111011110, 14'b11111111111010, 14'b00000000000000, 14'b11111111111101, 14'b00000000000011, 14'b11111111111111}, 
{14'b11111111101100, 14'b11111111110100, 14'b11111111110101, 14'b11111111100001, 14'b11111111110001, 14'b11111111111111, 14'b00000000001101, 14'b11111111110101, 14'b00000000011001, 14'b00000000000000, 14'b00000000000000, 14'b11111111111111, 14'b00000000011100, 14'b00000000000000, 14'b11111111111111, 14'b11111111110110, 14'b11111111111111, 14'b00000000000000, 14'b11111111111111, 14'b00000000000000, 14'b11111111111111, 14'b11111111111111, 14'b00000000000000, 14'b11111111111111, 14'b00000000000101, 14'b11111111101000, 14'b00000000000001, 14'b11111111111111, 14'b11111111110110, 14'b11111111111111, 14'b00000000000000, 14'b11111111111111}, 
{14'b11111111000010, 14'b11111111111000, 14'b11111111001111, 14'b00000000001111, 14'b00000000111110, 14'b11111111111111, 14'b11111111111100, 14'b00000000011110, 14'b11111111000111, 14'b11111111111010, 14'b00000000000000, 14'b11111111100110, 14'b11111111111111, 14'b00000000001001, 14'b11111111100111, 14'b00000001100000, 14'b11111111111110, 14'b00000000000101, 14'b00000000011010, 14'b00000000011111, 14'b00000000000000, 14'b11111111010101, 14'b00000000000000, 14'b00000000110100, 14'b11111111101000, 14'b00000001011001, 14'b11111111101100, 14'b11111111100101, 14'b11111111000011, 14'b11111111000100, 14'b00000000000000, 14'b00000000000110}, 
{14'b00000000000000, 14'b11111111111110, 14'b11111111110110, 14'b00000000000000, 14'b00000000100111, 14'b11111111111101, 14'b11111111110111, 14'b00000000001011, 14'b00000000001100, 14'b00000000000000, 14'b11111111111110, 14'b11111111111111, 14'b11111111111111, 14'b11111111110001, 14'b11111111111111, 14'b00000000000000, 14'b00000000000000, 14'b11111111111111, 14'b00000000000000, 14'b00000000001010, 14'b00000000000010, 14'b11111111111111, 14'b00000000000000, 14'b00000000000000, 14'b00000000000100, 14'b11111111101111, 14'b00000000001000, 14'b00000000011111, 14'b11111111111111, 14'b00000000000000, 14'b00000000000110, 14'b00000000001000}, 
{14'b00000000001100, 14'b00000000000000, 14'b11111111110010, 14'b11111111011111, 14'b11111110011010, 14'b00000000010001, 14'b00000000000000, 14'b11111110010110, 14'b00000000000100, 14'b11111111111111, 14'b00000000000000, 14'b11111111111111, 14'b00000000000001, 14'b00000000000000, 14'b11111111111101, 14'b11111111001111, 14'b11111111111111, 14'b00000000011100, 14'b00000000010000, 14'b00000000011000, 14'b11111111000111, 14'b11111111010010, 14'b00000000001111, 14'b11111111111011, 14'b11111111111010, 14'b00000000101101, 14'b11111111110011, 14'b11111111111111, 14'b11111111111111, 14'b00000000011011, 14'b11111111111111, 14'b00000000000000}, 
{14'b11111111100110, 14'b11111111000000, 14'b00000000000000, 14'b11111111111111, 14'b00000000101010, 14'b11111111011101, 14'b11111111100011, 14'b00000000001110, 14'b11111111111111, 14'b00000000010011, 14'b00000000001001, 14'b11111111110110, 14'b00000000000000, 14'b00000000000001, 14'b11111111111101, 14'b11111111011111, 14'b00000000010110, 14'b00000000000011, 14'b00000000100110, 14'b00000000001011, 14'b00000000000000, 14'b11111111111011, 14'b00000000010000, 14'b11111111110100, 14'b11111111011000, 14'b11111111111111, 14'b00000000010111, 14'b11111111111111, 14'b00000000000001, 14'b11111111110011, 14'b00000000010001, 14'b00000000100011}, 
{14'b00000000000001, 14'b00000000000000, 14'b00000000011100, 14'b00000000000001, 14'b11111111111010, 14'b00000000010111, 14'b00000000001011, 14'b11111111111111, 14'b00000000000000, 14'b11111111101110, 14'b11111111111001, 14'b11111111101010, 14'b11111111111111, 14'b00000000000110, 14'b11111111110111, 14'b00000001101011, 14'b00000000000000, 14'b11111111110011, 14'b11111111100111, 14'b11111111111110, 14'b00000000011001, 14'b00000000010000, 14'b00000000000000, 14'b11111111111111, 14'b00000000011100, 14'b00000000100010, 14'b00000000111111, 14'b00000000000001, 14'b00000000000000, 14'b00000000000000, 14'b11111111111110, 14'b11111111110110}, 
{14'b11111111101100, 14'b00000000000110, 14'b00000000000101, 14'b11111111100000, 14'b11111111011101, 14'b00000000111100, 14'b00000000000110, 14'b00000000000000, 14'b11111111101011, 14'b11111111110100, 14'b00000000010000, 14'b00000000001001, 14'b00000000000000, 14'b11111111110101, 14'b00000000100100, 14'b11111111111111, 14'b11111111111110, 14'b00000000000000, 14'b00000000000001, 14'b11111111111010, 14'b00000000001010, 14'b00000000000010, 14'b00000000001110, 14'b11111111111111, 14'b00000000000000, 14'b00000001010100, 14'b11111111111000, 14'b11111111111101, 14'b11111111111111, 14'b11111111110010, 14'b11111111111010, 14'b00000000010110}, 
{14'b00000000000111, 14'b00000000001001, 14'b00000000101001, 14'b11111111111010, 14'b00000000001100, 14'b00000000101100, 14'b00000000000000, 14'b11111111111100, 14'b00000000001111, 14'b11111111110001, 14'b11111111111111, 14'b11111111110000, 14'b00000000000000, 14'b00000000110010, 14'b11111111111101, 14'b00000000000000, 14'b00000000011110, 14'b00000000000000, 14'b00000000000000, 14'b11111111010111, 14'b11111111100000, 14'b11111111111011, 14'b11111111111111, 14'b11111111101101, 14'b11111111111011, 14'b11111111110101, 14'b11111111100110, 14'b11111111100100, 14'b00000000000011, 14'b00000000001110, 14'b11111111001101, 14'b00000000000000}, 
{14'b11111111011001, 14'b00000000000000, 14'b11111111111110, 14'b11111111111001, 14'b11111111111111, 14'b00000000010001, 14'b11111111110110, 14'b00000000100010, 14'b11111111010001, 14'b11111111111111, 14'b00000000000000, 14'b11111111111111, 14'b00000000000000, 14'b00000000000000, 14'b11111111111111, 14'b11111111110100, 14'b00000000001010, 14'b00000000010111, 14'b11111111111110, 14'b11111111011111, 14'b11111111111000, 14'b00000000001110, 14'b00000000001000, 14'b00000000000000, 14'b00000000000000, 14'b00000000001010, 14'b11111111100001, 14'b00000000000000, 14'b11111111111111, 14'b00000000000000, 14'b00000000000000, 14'b11111111101111}, 
{14'b11111111010100, 14'b11111111111111, 14'b11111111111111, 14'b11111111111101, 14'b11111111111111, 14'b00000000001101, 14'b00000000000000, 14'b00000000000100, 14'b00000000000100, 14'b00000000001000, 14'b00000000001010, 14'b00000000010100, 14'b00000000000011, 14'b11111111110011, 14'b00000000000000, 14'b00000000110000, 14'b00000000000000, 14'b00000000000000, 14'b11111111111111, 14'b00000000001110, 14'b00000000010010, 14'b00000000000011, 14'b00000000000101, 14'b11111111111100, 14'b11111111111011, 14'b00000000000011, 14'b11111111110111, 14'b11111111101111, 14'b00000000011010, 14'b11111111111100, 14'b00000000000100, 14'b11111111100111}, 
{14'b00000000000000, 14'b11111111111111, 14'b00000000000100, 14'b00000000000000, 14'b00000001110100, 14'b11111111111111, 14'b00000000000000, 14'b11111111111111, 14'b00000000001110, 14'b11111111110110, 14'b00000000000000, 14'b00000000000000, 14'b00000000000000, 14'b00000000010000, 14'b00000000000000, 14'b11111111101101, 14'b11111111111111, 14'b11111111110111, 14'b00000000101001, 14'b00000000000000, 14'b11111111111111, 14'b11111111111111, 14'b00000000000000, 14'b11111111111111, 14'b00000000000000, 14'b00000000001000, 14'b00000000000000, 14'b00000000000000, 14'b11111111111111, 14'b11111111111111, 14'b00000000000000, 14'b00000000000101}, 
{14'b11111111111111, 14'b00000000000011, 14'b11111111111111, 14'b00000000000110, 14'b11111111111010, 14'b11111111110000, 14'b11111111111000, 14'b00000000100011, 14'b00000000000000, 14'b00000000001100, 14'b11111111111110, 14'b00000000001000, 14'b11111111111011, 14'b11111111101011, 14'b11111111100111, 14'b00000000000001, 14'b11111111111111, 14'b11111111111011, 14'b00000000000000, 14'b00000000000000, 14'b11111111111111, 14'b00000000001001, 14'b00000000000100, 14'b11111111101111, 14'b00000000001110, 14'b11111111101010, 14'b00000000000000, 14'b00000000000000, 14'b11111111101010, 14'b00000000000000, 14'b00000000000101, 14'b11111111111100}, 
{14'b11111111111110, 14'b11111111110011, 14'b00000000000000, 14'b11111111111000, 14'b00000000011011, 14'b11111111111111, 14'b11111111111101, 14'b00000000001101, 14'b11111111001101, 14'b00000000000000, 14'b11111111111011, 14'b11111111111111, 14'b00000000101100, 14'b00000000011101, 14'b11111111110011, 14'b11111111111101, 14'b11111111111111, 14'b00000000000000, 14'b11111111111111, 14'b00000000000000, 14'b00000000000000, 14'b11111111101110, 14'b11111111110000, 14'b00000000010000, 14'b00000000000000, 14'b11111111101110, 14'b00000000000011, 14'b11111111110101, 14'b11111111111011, 14'b00000000010001, 14'b00000000000000, 14'b11111111100000}, 
{14'b00000001010001, 14'b00000000101011, 14'b11111111100000, 14'b00000000000000, 14'b11111111010011, 14'b00000000000000, 14'b00000000011100, 14'b00000000000011, 14'b00000000011100, 14'b11111111111111, 14'b11111111101100, 14'b11111111110101, 14'b00000000010010, 14'b00000000000011, 14'b11111111110011, 14'b00000000010000, 14'b00000001000100, 14'b11111111101111, 14'b11111111011010, 14'b00000000000000, 14'b11111111111100, 14'b11111111101001, 14'b11111111111110, 14'b11111111111111, 14'b00000000001011, 14'b11111111010001, 14'b00000000001011, 14'b11111111111111, 14'b00000000000000, 14'b00000000001101, 14'b11111111111100, 14'b00000000000111}, 
{14'b11111111110100, 14'b11111111100111, 14'b11111111111011, 14'b11111111101010, 14'b11111111111101, 14'b00000000000110, 14'b00000000000000, 14'b11111111111110, 14'b00000000000100, 14'b11111111111111, 14'b00000000000000, 14'b11111111100100, 14'b00000000001101, 14'b00000000001010, 14'b11111111110010, 14'b00000000111000, 14'b11111111111111, 14'b00000000000000, 14'b11111111111111, 14'b00000000000000, 14'b00000000101000, 14'b11111111000011, 14'b11111111110010, 14'b11111111111000, 14'b11111111111101, 14'b00000000011001, 14'b11111111111001, 14'b00000000000010, 14'b00000000111101, 14'b11111110111110, 14'b11111111010001, 14'b00000000000010}, 
{14'b00000000000010, 14'b11111111111000, 14'b11111111111111, 14'b00000000000000, 14'b11111110100011, 14'b11111110110010, 14'b00000000000000, 14'b11111111111111, 14'b11111111011110, 14'b00000000000011, 14'b00000000000000, 14'b11111111111100, 14'b00000000000000, 14'b11111111111000, 14'b11111111111001, 14'b11111111110111, 14'b11111111101101, 14'b00000000100100, 14'b00000000000000, 14'b00000000000101, 14'b11111111111111, 14'b11111111110110, 14'b00000000000000, 14'b11111111110100, 14'b00000000011100, 14'b11111110110000, 14'b00000000011100, 14'b11111111111111, 14'b11111111111111, 14'b00000000011001, 14'b11111111111111, 14'b00000000011110}, 
{14'b11111111111111, 14'b00000000000000, 14'b11111111111010, 14'b00000000001001, 14'b00000000000111, 14'b11111111010100, 14'b00000000000000, 14'b00000000001000, 14'b00000001001010, 14'b11111111111110, 14'b00000000000000, 14'b00000000000111, 14'b00000000101101, 14'b11111111111011, 14'b00000000000001, 14'b00000000001100, 14'b11111111111111, 14'b00000000000011, 14'b11111111111111, 14'b00000000000000, 14'b11111111011100, 14'b00000000000100, 14'b00000000001000, 14'b00000000000010, 14'b11111111111111, 14'b00000000011011, 14'b00000000000000, 14'b00000000010000, 14'b11111111001010, 14'b00000000001101, 14'b00000000110010, 14'b00000000000000}, 
{14'b11111111010011, 14'b00000000011011, 14'b11111111011110, 14'b00000000001111, 14'b11111111110010, 14'b00000000000000, 14'b00000000111111, 14'b11111111100010, 14'b11111111011010, 14'b00000000010101, 14'b11111111100011, 14'b11111111111100, 14'b11111111111111, 14'b00000000101100, 14'b11111111111111, 14'b11111111011001, 14'b11111111111111, 14'b00000000111000, 14'b11111111000011, 14'b11111111111100, 14'b00000000101000, 14'b11111111010001, 14'b00000000000110, 14'b11111111111110, 14'b00000000100010, 14'b11111110111110, 14'b11111111010001, 14'b11111111100110, 14'b11111111111111, 14'b00000000001101, 14'b00000000000011, 14'b00000000010110}, 
{14'b11111111110100, 14'b00000000000110, 14'b11111111111111, 14'b00000000010011, 14'b11111111111011, 14'b00000000011101, 14'b00000000000000, 14'b11111111111110, 14'b11111111111111, 14'b00000000000000, 14'b00000000000000, 14'b11111111111111, 14'b11111111111111, 14'b00000001000010, 14'b00000000000001, 14'b00000000011000, 14'b00000000000000, 14'b11111111100100, 14'b11111111110110, 14'b11111111111111, 14'b11111111111101, 14'b00000000000101, 14'b11111111111111, 14'b11111111101000, 14'b11111111111111, 14'b00000000100101, 14'b00000000100111, 14'b11111111111111, 14'b11111111111101, 14'b00000000000000, 14'b11111111111111, 14'b11111111110011}, 
{14'b11111111110101, 14'b00000000000000, 14'b00000000100010, 14'b00000000000000, 14'b00000000000000, 14'b11111111110001, 14'b00000000000000, 14'b11111110010001, 14'b00000000011011, 14'b00000000000001, 14'b00000000000011, 14'b11111111010001, 14'b00000000000000, 14'b11111111101110, 14'b11111111111011, 14'b00000000000000, 14'b00000000000010, 14'b00000000000000, 14'b00000000001110, 14'b00000000000000, 14'b11111111111110, 14'b00000000101010, 14'b00000000110000, 14'b11111111100011, 14'b11111111101101, 14'b00000000011111, 14'b11111111011000, 14'b00000000000011, 14'b11111111111111, 14'b11111111111111, 14'b11111111111111, 14'b00000000010111}, 
{14'b11111111110001, 14'b11111111111111, 14'b11111111100001, 14'b11111111100110, 14'b11111111111110, 14'b11111111101110, 14'b00000000000000, 14'b00000000001011, 14'b11111111100001, 14'b11111111110101, 14'b11111111111001, 14'b00000000000000, 14'b00000000000011, 14'b11111111111110, 14'b11111111111000, 14'b00000000001100, 14'b00000000011100, 14'b00000000010000, 14'b11111111101111, 14'b00000000000110, 14'b11111111111110, 14'b11111111111100, 14'b00000000000010, 14'b00000000000010, 14'b11111111110111, 14'b00000000001011, 14'b11111111110100, 14'b00000000000111, 14'b11111111111111, 14'b11111111011010, 14'b11111111111100, 14'b00000000011100}, 
{14'b11111111111100, 14'b11111111110101, 14'b00000000001001, 14'b00000000100000, 14'b00000000001010, 14'b00000000001010, 14'b00000000000101, 14'b11111111100110, 14'b11111111100101, 14'b00000000001000, 14'b00000000000001, 14'b00000000000101, 14'b00000000000010, 14'b00000000000000, 14'b00000000011010, 14'b00000000000000, 14'b11111111111001, 14'b00000000001101, 14'b11111111111100, 14'b11111111111011, 14'b00000000001110, 14'b11111111110000, 14'b11111111111100, 14'b00000000010000, 14'b00000000000010, 14'b11111111110010, 14'b11111111100110, 14'b11111111111110, 14'b11111111011100, 14'b00000000000111, 14'b00000000001101, 14'b00000000000000}, 
{14'b11111111111110, 14'b11111111111101, 14'b11111111111110, 14'b11111111111011, 14'b11111111101111, 14'b11111111101110, 14'b00000000001000, 14'b00000000000001, 14'b11111111101000, 14'b00000000010101, 14'b11111111111101, 14'b11111111111111, 14'b11111111110001, 14'b00000000000000, 14'b00000000000011, 14'b11111111111001, 14'b11111111111101, 14'b11111111111010, 14'b11111111110101, 14'b00000000000000, 14'b11111111101110, 14'b00000000001101, 14'b11111111100100, 14'b00000000000000, 14'b00000000000101, 14'b00000000001111, 14'b00000000000011, 14'b00000000000000, 14'b00000000100101, 14'b00000000000110, 14'b00000000000000, 14'b00000000001010}, 
{14'b11111111111101, 14'b00000000100000, 14'b11111111111111, 14'b11111111111011, 14'b11111111100100, 14'b11111111110110, 14'b00000000110100, 14'b11111110100111, 14'b11111111010011, 14'b11111111100110, 14'b11111111100011, 14'b11111111011111, 14'b11111111111111, 14'b00000000111101, 14'b11111111111100, 14'b00000000000000, 14'b11111111100100, 14'b00000000111001, 14'b11111111001011, 14'b00000000000000, 14'b11111111111111, 14'b11111111010100, 14'b00000000000000, 14'b11111111111111, 14'b00000000000111, 14'b11111111111000, 14'b11111111101101, 14'b11111111111111, 14'b00000000010110, 14'b00000000000000, 14'b11111111110101, 14'b00000000000000}, 
{14'b00000000101111, 14'b11111111110001, 14'b00000000010000, 14'b11111111111011, 14'b00000000001001, 14'b11111111111111, 14'b11111111111111, 14'b11111111110100, 14'b00000000000000, 14'b00000000001011, 14'b11111111111111, 14'b11111111111000, 14'b11111111111111, 14'b00000000011101, 14'b00000000000010, 14'b00000000000101, 14'b00000000000011, 14'b11111111111100, 14'b00000000000010, 14'b00000000000000, 14'b11111111111110, 14'b11111111111111, 14'b11111111011000, 14'b11111111111111, 14'b00000000000111, 14'b11111111110001, 14'b11111111101110, 14'b11111111111111, 14'b11111111111111, 14'b00000001000111, 14'b11111111011011, 14'b11111111110001}, 
{14'b11111111111010, 14'b11111111110010, 14'b11111111110111, 14'b00000000000100, 14'b00000000010001, 14'b11111111101111, 14'b11111111111111, 14'b11111111100011, 14'b00000000000111, 14'b00000000010001, 14'b11111111100100, 14'b11111111011111, 14'b00000000000011, 14'b11111110101000, 14'b11111111110110, 14'b11111111110000, 14'b11111111100110, 14'b11111111111111, 14'b00000000010001, 14'b00000000000000, 14'b11111111111010, 14'b11111111111010, 14'b00000000000000, 14'b00000000000000, 14'b11111111111000, 14'b11111110011111, 14'b11111110111000, 14'b11111111011101, 14'b00000000000111, 14'b00000000011010, 14'b11111111111111, 14'b00000000011110}, 
{14'b11111111110100, 14'b11111111100100, 14'b00000000010100, 14'b00000000001001, 14'b00000000000101, 14'b11111111110100, 14'b11111111111011, 14'b00000000001100, 14'b00000001000100, 14'b11111111101010, 14'b11111111111111, 14'b11111111111111, 14'b00000000001111, 14'b11111111111000, 14'b11111111111101, 14'b11111111111101, 14'b11111111110011, 14'b11111111111111, 14'b00000000000000, 14'b00000000011101, 14'b11111111101110, 14'b11111111111111, 14'b00000000010000, 14'b11111111111110, 14'b00000000000000, 14'b00000001000011, 14'b00000000101001, 14'b00000000000000, 14'b00000000000000, 14'b11111111001010, 14'b11111111110111, 14'b11111111111111}, 
{14'b00000000000001, 14'b00000000000110, 14'b11111111111110, 14'b00000000000000, 14'b00000000011101, 14'b11111111000010, 14'b00000000000000, 14'b11111111110011, 14'b00000000010111, 14'b00000000000000, 14'b11111111111101, 14'b00000000000000, 14'b00000000000000, 14'b11111111111111, 14'b00000000000000, 14'b11111111110010, 14'b00000000100001, 14'b11111111111111, 14'b11111111111110, 14'b11111111111111, 14'b00000000000000, 14'b11111111111111, 14'b00000000000000, 14'b11111111111111, 14'b00000000000001, 14'b11111111010111, 14'b00000000000110, 14'b00000000010111, 14'b11111111111111, 14'b00000000001100, 14'b11111111111111, 14'b00000000001001}, 
{14'b11111111100110, 14'b00000000000001, 14'b11111111000010, 14'b00000000000000, 14'b11111111111001, 14'b11111111111010, 14'b11111111111111, 14'b11111111110100, 14'b11111111111011, 14'b11111111110111, 14'b00000000000110, 14'b00000000000011, 14'b11111111101001, 14'b00000000000000, 14'b11111111111111, 14'b11111111111110, 14'b00000000001001, 14'b11111111111101, 14'b11111111111100, 14'b11111111111100, 14'b11111111111111, 14'b00000000100010, 14'b11111111111111, 14'b00000000000000, 14'b11111111111110, 14'b00000000101000, 14'b00000000011000, 14'b00000000000100, 14'b11111111110011, 14'b11111111111110, 14'b00000000001000, 14'b00000000000111}, 
{14'b00000000000100, 14'b00000000000101, 14'b11111111111111, 14'b00000000000000, 14'b11111111000100, 14'b00000000000101, 14'b00000000000011, 14'b11111111111111, 14'b00000000000000, 14'b11111111101010, 14'b11111111111111, 14'b00000000000000, 14'b11111111101011, 14'b00000000000000, 14'b00000000000000, 14'b00000000000000, 14'b00000000000000, 14'b11111111010010, 14'b00000000000001, 14'b11111111111111, 14'b11111111111111, 14'b00000000000000, 14'b00000000010000, 14'b11111111111111, 14'b00000000000000, 14'b00000000111010, 14'b00000000101011, 14'b00000000000000, 14'b00000000000000, 14'b11111111100010, 14'b00000000000000, 14'b11111111111111}, 
{14'b00000000001001, 14'b00000000000110, 14'b00000000100000, 14'b11111111100000, 14'b00000000010000, 14'b00000000001111, 14'b00000000000000, 14'b00000000011000, 14'b00000000000001, 14'b11111111111110, 14'b00000000000100, 14'b00000000000000, 14'b11111111111111, 14'b00000000001111, 14'b11111111111111, 14'b11111111111010, 14'b00000000000000, 14'b00000000000100, 14'b11111111111001, 14'b00000000001100, 14'b00000000000100, 14'b11111110110101, 14'b11111111110001, 14'b00000000001011, 14'b11111111111111, 14'b11111110111111, 14'b11111111101111, 14'b11111111111101, 14'b11111111111111, 14'b11111111111000, 14'b00000000000000, 14'b11111111111010}, 
{14'b00000000000000, 14'b11111111111111, 14'b11111111110100, 14'b11111111101010, 14'b00000000000101, 14'b00000000000000, 14'b00000000001100, 14'b11111111111111, 14'b00000000011111, 14'b11111111111111, 14'b00000000000000, 14'b11111111010100, 14'b11111111111111, 14'b00000000010000, 14'b11111111111111, 14'b11111111011110, 14'b00000000000000, 14'b11111111111110, 14'b00000000100001, 14'b11111111111111, 14'b11111111001000, 14'b11111111111111, 14'b00000000100001, 14'b11111111111111, 14'b11111111111111, 14'b00000000010001, 14'b11111111110011, 14'b00000000001000, 14'b00000000000000, 14'b11111111100110, 14'b00000000000000, 14'b00000000000000}, 
{14'b11111111100100, 14'b00000000000000, 14'b00000000000000, 14'b11111111111111, 14'b00000000111111, 14'b11111111110000, 14'b11111111111111, 14'b11111111111111, 14'b11111111111010, 14'b11111111111001, 14'b00000000001000, 14'b00000000010001, 14'b11111111111011, 14'b00000000011111, 14'b00000000000000, 14'b11111111111111, 14'b11111111011011, 14'b11111111111111, 14'b00000000000000, 14'b11111111110101, 14'b00000000000000, 14'b00000000000100, 14'b00000000000001, 14'b11111111111110, 14'b11111111111001, 14'b11111111100110, 14'b11111111011010, 14'b00000000000000, 14'b11111111110001, 14'b00000000000101, 14'b11111111111111, 14'b00000000001001}, 
{14'b11111111001011, 14'b11111111101011, 14'b11111111101100, 14'b00000000000000, 14'b00000001001001, 14'b11111111100011, 14'b00000000000000, 14'b11111111111001, 14'b11111111001011, 14'b00000000010001, 14'b11111111111111, 14'b00000001001000, 14'b00000000000000, 14'b11111111111001, 14'b11111111111111, 14'b00000000000100, 14'b11111111111101, 14'b00000000000000, 14'b11111111111010, 14'b00000000111111, 14'b00000000000100, 14'b11111111111010, 14'b00000000001110, 14'b11111111111111, 14'b11111111111111, 14'b11111111110011, 14'b11111111111010, 14'b11111111000100, 14'b11111111101101, 14'b11111111111111, 14'b11111111111111, 14'b11111111111000}, 
{14'b00000000011100, 14'b11111110011001, 14'b11111110100011, 14'b11111111101010, 14'b00000001010101, 14'b11111111111111, 14'b11111111010011, 14'b00000000100001, 14'b00000000000111, 14'b00000000000000, 14'b00000000011010, 14'b11111111011101, 14'b00000000000000, 14'b00000000000000, 14'b11111111111011, 14'b00000000000010, 14'b11111111110010, 14'b11111110001010, 14'b00000000010101, 14'b00000000101100, 14'b00000000100001, 14'b00000000000000, 14'b00000000000011, 14'b11111111001100, 14'b11111110101111, 14'b11111111111111, 14'b11111111011001, 14'b11111111000101, 14'b11111111100111, 14'b11111110001111, 14'b00000000110101, 14'b00000000110110}, 
{14'b00000000000000, 14'b00000000000000, 14'b00000000000000, 14'b00000000000000, 14'b00000000100001, 14'b11111111101000, 14'b00000000000010, 14'b00000000001001, 14'b11111111010011, 14'b00000000000100, 14'b11111111111111, 14'b11111111111111, 14'b11111111111111, 14'b00000000011110, 14'b00000000000110, 14'b00000000000010, 14'b00000000000111, 14'b00000000101010, 14'b11111111100100, 14'b00000000000000, 14'b11111111101010, 14'b11111111111111, 14'b00000000101000, 14'b00000000000001, 14'b11111111111111, 14'b11111110111000, 14'b11111111111110, 14'b11111111101100, 14'b11111111111000, 14'b00000000000000, 14'b00000000010001, 14'b00000000001101}, 
{14'b11111111111010, 14'b00000000010001, 14'b11111111011001, 14'b00000000000010, 14'b00000000011000, 14'b11111111111010, 14'b11111111111111, 14'b00000000010100, 14'b00000000000000, 14'b11111111111111, 14'b11111111110111, 14'b00000000000000, 14'b00000000000000, 14'b11111111111011, 14'b11111111110000, 14'b11111111110111, 14'b11111111111000, 14'b11111111110111, 14'b11111111110001, 14'b00000000000000, 14'b11111111111111, 14'b11111111111010, 14'b11111111110111, 14'b00000000110010, 14'b00000000000000, 14'b11111111010001, 14'b11111111111110, 14'b00000000001111, 14'b00000000000000, 14'b00000000000000, 14'b00000000100000, 14'b11111111111111}, 
{14'b11111111111111, 14'b00000000000000, 14'b11111111111111, 14'b11111111101100, 14'b11111110010001, 14'b00000000000000, 14'b00000000000000, 14'b11111111111111, 14'b11111110110011, 14'b00000000001010, 14'b11111111110011, 14'b11111111111111, 14'b00000000000000, 14'b11111111010000, 14'b11111111111010, 14'b11111111111111, 14'b00000000000000, 14'b00000000000001, 14'b00000000000100, 14'b00000000101100, 14'b11111111110000, 14'b11111111011001, 14'b00000000000000, 14'b11111111011110, 14'b11111111110011, 14'b11111111100010, 14'b11111111111111, 14'b11111111111110, 14'b11111111111101, 14'b11111111000011, 14'b11111111111011, 14'b00000000011111}, 
{14'b00000000001110, 14'b00000000011100, 14'b11111111111111, 14'b00000000010100, 14'b11111111100101, 14'b11111111110000, 14'b00000000001100, 14'b00000000001000, 14'b11111111111001, 14'b11111111111111, 14'b11111111111111, 14'b11111111111111, 14'b11111111111111, 14'b11111111010110, 14'b11111111111111, 14'b00000000010010, 14'b11111111110001, 14'b00000000000100, 14'b11111111111111, 14'b11111111111111, 14'b00000000011010, 14'b11111111010110, 14'b00000000100011, 14'b00000000000110, 14'b00000000000000, 14'b00000000011011, 14'b00000000000000, 14'b11111111111011, 14'b11111111001111, 14'b11111111110001, 14'b11111111101010, 14'b00000000010110}, 
{14'b00000000000000, 14'b00000000000000, 14'b11111111010001, 14'b11111111111111, 14'b00000000011010, 14'b11111111101101, 14'b11111111111110, 14'b11111111111111, 14'b00000000000010, 14'b00000000000000, 14'b00000000000000, 14'b11111111100101, 14'b00000000001100, 14'b00000000000000, 14'b00000000000000, 14'b00000000000100, 14'b11111111111111, 14'b11111111101100, 14'b00000000000010, 14'b00000000000000, 14'b11111111111011, 14'b11111111111101, 14'b00000000100101, 14'b11111111111111, 14'b00000000000000, 14'b11111111011010, 14'b11111111010110, 14'b00000000011110, 14'b11111111111111, 14'b11111111111111, 14'b00000000000011, 14'b00000000100100}, 
{14'b11111111010100, 14'b11111111111111, 14'b11111111100100, 14'b00000000000000, 14'b11111111010010, 14'b00000000000000, 14'b11111111111111, 14'b11111111110111, 14'b11111110111011, 14'b11111111111100, 14'b00000000000000, 14'b11111111111110, 14'b11111111111111, 14'b00000000000000, 14'b11111111111110, 14'b11111111111001, 14'b11111111101101, 14'b11111111110011, 14'b00000000001000, 14'b11111111111111, 14'b11111111111100, 14'b00000000000000, 14'b00000000101011, 14'b11111111111111, 14'b00000000010011, 14'b00000000001011, 14'b11111111101110, 14'b00000000011011, 14'b11111111111010, 14'b00000000000000, 14'b11111111111111, 14'b00000001001010}, 
{14'b11111111010111, 14'b00000000000011, 14'b00000000000110, 14'b11111111111100, 14'b00000000011111, 14'b11111111011001, 14'b11111111111111, 14'b00000000100001, 14'b00000000010100, 14'b00000000000001, 14'b11111111111111, 14'b11111111110111, 14'b11111111110100, 14'b11111111110111, 14'b11111111111001, 14'b00000000001011, 14'b11111111111111, 14'b00000000000001, 14'b00000000010010, 14'b00000000000000, 14'b00000000000000, 14'b00000000000001, 14'b00000000100000, 14'b00000000000101, 14'b00000000000000, 14'b11111111110010, 14'b11111111111111, 14'b00000000000000, 14'b11111111111110, 14'b11111111111110, 14'b11111111111111, 14'b00000000001000}, 
{14'b11111111111111, 14'b00000000000000, 14'b11111111100100, 14'b11111111110110, 14'b00000000100100, 14'b11111111111111, 14'b11111111110110, 14'b00000000011111, 14'b11111111111001, 14'b00000000100101, 14'b00000000001010, 14'b11111111110000, 14'b00000000000000, 14'b00000000000000, 14'b11111111111110, 14'b00000000000010, 14'b11111111110110, 14'b11111111011110, 14'b00000000100011, 14'b00000000010011, 14'b00000001010001, 14'b00000000011001, 14'b00000000011111, 14'b11111111111111, 14'b00000000000000, 14'b00000000000000, 14'b00000000000111, 14'b00000000001010, 14'b11111111001010, 14'b11111111111111, 14'b11111111111111, 14'b11111111111111}, 
{14'b00000000000000, 14'b11111111110100, 14'b11111111110010, 14'b00000000000000, 14'b11111111100000, 14'b00000000000000, 14'b00000000011000, 14'b00000000001101, 14'b00000000000110, 14'b11111111110011, 14'b00000000000000, 14'b11111111111111, 14'b11111111111111, 14'b11111111111111, 14'b11111111111010, 14'b00000000011001, 14'b11111111111111, 14'b11111111111111, 14'b11111111011001, 14'b00000000000000, 14'b11111111100111, 14'b11111111111111, 14'b00000000000000, 14'b11111111111111, 14'b00000000000001, 14'b00000000000010, 14'b00000000000011, 14'b00000000010001, 14'b11111111110111, 14'b11111111111111, 14'b11111111000110, 14'b00000000001010}, 
{14'b00000000111000, 14'b11111111111110, 14'b00000000001000, 14'b11111111110010, 14'b11111111110101, 14'b00000000000100, 14'b00000000010100, 14'b00000000000000, 14'b00000001000011, 14'b00000000000000, 14'b11111111111101, 14'b00000000000010, 14'b00000000001100, 14'b11111111111111, 14'b00000000000110, 14'b00000000001101, 14'b11111111111111, 14'b11111111000111, 14'b11111111111000, 14'b11111111111111, 14'b00000000001110, 14'b00000000000000, 14'b11111111111111, 14'b00000000001110, 14'b00000000000010, 14'b11111111011110, 14'b11111111110010, 14'b00000000010000, 14'b11111111111100, 14'b00000000100001, 14'b11111111111111, 14'b11111111101001}, 
{14'b00000000000001, 14'b00000000001101, 14'b11111111111111, 14'b11111111111011, 14'b11111111010010, 14'b11111111111111, 14'b00000000000101, 14'b11111111111010, 14'b00000000010101, 14'b11111111111011, 14'b11111111111111, 14'b11111111111011, 14'b11111111111111, 14'b11111111111011, 14'b00000000000000, 14'b00000000101000, 14'b00000000000000, 14'b11111111111111, 14'b11111111111111, 14'b11111111111111, 14'b11111111111111, 14'b11111111111111, 14'b00000000000100, 14'b00000000010000, 14'b00000000000000, 14'b00000000000000, 14'b00000000000100, 14'b11111111111111, 14'b00000000000000, 14'b00000000000010, 14'b00000000000000, 14'b00000000001100}, 
{14'b11111111011000, 14'b00000000010000, 14'b00000000000010, 14'b11111111110010, 14'b11111111001100, 14'b11111111111101, 14'b00000000001000, 14'b11111111001101, 14'b00000001000001, 14'b00000000001001, 14'b00000000000010, 14'b00000000001100, 14'b00000000000101, 14'b00000000000000, 14'b00000000110100, 14'b11111111110101, 14'b00000000000000, 14'b00000000000000, 14'b11111111111111, 14'b00000000000000, 14'b11111111001000, 14'b00000000000010, 14'b00000000010011, 14'b00000000000100, 14'b00000000000100, 14'b11111110101011, 14'b11111111010100, 14'b11111111100001, 14'b00000000000000, 14'b11111111111111, 14'b00000000101001, 14'b11111111100101}, 
{14'b11111111111110, 14'b11111111100111, 14'b11111111110010, 14'b11111111001011, 14'b11111111011110, 14'b00000000101011, 14'b00000000100111, 14'b11111111101010, 14'b00000000000101, 14'b11111111111011, 14'b11111111110011, 14'b11111111011111, 14'b00000000001101, 14'b11111111011011, 14'b00000000011000, 14'b11111111111111, 14'b00000000101010, 14'b11111111111111, 14'b11111111111111, 14'b11111111101110, 14'b11111111111010, 14'b11111111110111, 14'b11111111011101, 14'b00000000001010, 14'b11111111111111, 14'b11111111111111, 14'b11111111100010, 14'b00000000101000, 14'b00000000100011, 14'b11111111110100, 14'b11111110101111, 14'b00000000010010}, 
{14'b00000000000000, 14'b11111111111100, 14'b11111111111111, 14'b11111111110011, 14'b00000000000011, 14'b00000000000001, 14'b00000000001000, 14'b00000000000000, 14'b00000000001111, 14'b11111111111111, 14'b00000000000000, 14'b00000000001100, 14'b00000000000000, 14'b00000000000001, 14'b11111111101111, 14'b11111111110010, 14'b00000000000000, 14'b00000000010111, 14'b00000000000111, 14'b00000000010000, 14'b11111111111101, 14'b11111111101011, 14'b11111111111111, 14'b00000000001001, 14'b11111111111111, 14'b00000000000100, 14'b11111111111111, 14'b00000000001000, 14'b00000000000000, 14'b00000000001010, 14'b11111111001111, 14'b11111111111111}, 
{14'b00000000100111, 14'b11111111111110, 14'b00000000010011, 14'b11111111011000, 14'b11111111100111, 14'b11111111111111, 14'b11111111111111, 14'b00000000000011, 14'b00000000000000, 14'b11111111101111, 14'b00000000000000, 14'b00000000000000, 14'b00000000000000, 14'b00000000000000, 14'b11111111101111, 14'b00000000010010, 14'b11111111111111, 14'b11111111111100, 14'b00000000000000, 14'b00000000001111, 14'b11111111100110, 14'b00000000001110, 14'b00000000010001, 14'b00000000010000, 14'b11111111111111, 14'b00000001000110, 14'b11111111101100, 14'b00000000101110, 14'b11111111111001, 14'b11111111010001, 14'b11111111101001, 14'b00000000010001}, 
{14'b11111110111010, 14'b11111111111100, 14'b11111111101100, 14'b11111111111111, 14'b00000000100001, 14'b11111111101001, 14'b11111111111000, 14'b00000000011110, 14'b00000000001100, 14'b11111111100001, 14'b00000000000000, 14'b11111111111100, 14'b11111111111110, 14'b00000000010001, 14'b11111111100000, 14'b11111111111110, 14'b00000000000000, 14'b11111111111111, 14'b11111111111101, 14'b00000000000000, 14'b11111111100111, 14'b11111111111111, 14'b00000000000000, 14'b11111111010101, 14'b00000000001000, 14'b00000001001111, 14'b00000000101100, 14'b11111111111011, 14'b11111111101011, 14'b11111111000110, 14'b00000000000000, 14'b11111111111001}, 
{14'b00000000000010, 14'b00000000011011, 14'b00000000000010, 14'b11111111101100, 14'b00000000000000, 14'b11111111111100, 14'b00000000000000, 14'b00000000011010, 14'b00000000011011, 14'b11111111101110, 14'b00000000010001, 14'b00000000000011, 14'b11111111111111, 14'b11111111111110, 14'b11111111101011, 14'b00000000100000, 14'b11111111111010, 14'b11111111010110, 14'b00000000001110, 14'b11111111111111, 14'b11111111111111, 14'b00000000001110, 14'b11111111110110, 14'b11111111111111, 14'b11111111111001, 14'b00000000001011, 14'b11111111101110, 14'b00000000010001, 14'b11111111010001, 14'b00000000001010, 14'b11111111111111, 14'b00000000010100}, 
{14'b11111111111010, 14'b00000000000000, 14'b00000000001011, 14'b00000000000000, 14'b11111111111000, 14'b11111111111111, 14'b00000000001101, 14'b11111111111111, 14'b00000000000000, 14'b00000000000000, 14'b00000000000000, 14'b00000000000010, 14'b11111111110010, 14'b00000000000001, 14'b00000000001110, 14'b00000000000101, 14'b00000000001101, 14'b11111111111111, 14'b11111111111111, 14'b00000000010000, 14'b00000000011111, 14'b11111111110011, 14'b00000000000000, 14'b11111111111111, 14'b00000000000001, 14'b11111111000100, 14'b11111111111111, 14'b11111111110110, 14'b11111111111111, 14'b00000001001000, 14'b00000000000000, 14'b11111111100101}, 
{14'b11111111111100, 14'b11111111110000, 14'b11111111111110, 14'b00000000000000, 14'b00000000001011, 14'b11111111111111, 14'b00000000000000, 14'b11111111111101, 14'b00000000001001, 14'b11111111111110, 14'b00000000000000, 14'b00000000000100, 14'b00000000100101, 14'b11111111110010, 14'b00000000000001, 14'b11111110010011, 14'b11111111111110, 14'b11111111111000, 14'b00000000000001, 14'b11111111111001, 14'b00000000001011, 14'b11111111100011, 14'b00000000001110, 14'b00000000001101, 14'b11111111111110, 14'b11111110100100, 14'b11111111100010, 14'b11111111111101, 14'b11111111111101, 14'b00000000110001, 14'b11111111111111, 14'b00000000010011}, 
{14'b00000000000110, 14'b00000000000000, 14'b00000000010110, 14'b11111111110001, 14'b11111111110111, 14'b00000000011110, 14'b11111111101011, 14'b00000000000111, 14'b11111111011000, 14'b00000000000001, 14'b00000000000010, 14'b11111111110101, 14'b00000000000000, 14'b00000000000000, 14'b11111111100111, 14'b00000000110111, 14'b11111111100000, 14'b11111111111110, 14'b00000000001111, 14'b11111111111111, 14'b00000000001000, 14'b11111111000010, 14'b00000000101000, 14'b11111111111111, 14'b11111111110000, 14'b00000000111110, 14'b00000000010010, 14'b11111111101011, 14'b11111111101110, 14'b11111110111011, 14'b11111111111110, 14'b00000000000010}, 
{14'b11111111111111, 14'b00000000000000, 14'b11111111111011, 14'b11111111011101, 14'b11111111111111, 14'b11111111001101, 14'b00000000000000, 14'b00000000100110, 14'b00000000011111, 14'b00000000000010, 14'b00000000000000, 14'b11111111110001, 14'b00000000101010, 14'b11111111111111, 14'b11111111111111, 14'b11111111111111, 14'b00000000110111, 14'b00000000000000, 14'b11111111111010, 14'b11111111111001, 14'b11111111010110, 14'b00000000010000, 14'b00000000000000, 14'b00000000000000, 14'b00000000000100, 14'b11111111110110, 14'b11111111000101, 14'b00000000100011, 14'b11111111000111, 14'b00000000000110, 14'b11111111110101, 14'b00000000000000}, 
{14'b00000000000111, 14'b00000000010111, 14'b00000000000001, 14'b11111111111111, 14'b11111111000101, 14'b00000000000000, 14'b11111111111111, 14'b00000000011111, 14'b00000000100011, 14'b11111111111111, 14'b11111111111111, 14'b11111111111111, 14'b00000000000000, 14'b00000000000000, 14'b00000000000000, 14'b00000000000000, 14'b00000000000000, 14'b11111111111111, 14'b00000000010101, 14'b11111111110010, 14'b11111111001000, 14'b11111111111011, 14'b11111111110011, 14'b11111111110011, 14'b11111111110111, 14'b11111111111111, 14'b11111111110111, 14'b11111111111101, 14'b11111111111110, 14'b00000000010010, 14'b11111111111111, 14'b00000000111011}
};

localparam logic signed [13:0] bias [32] = '{
14'b00000010111100,  // 1.474280834197998
14'b00000001011000,  // 0.6914801001548767
14'b00000010111000,  // 1.4406442642211914
14'b00000010110100,  // 1.408045768737793
14'b00000001111110,  // 0.9864811301231384
14'b00000001101110,  // 0.8636202812194824
14'b11111110110001,  // -0.6153604388237
14'b00000000111101,  // 0.4839226007461548
14'b00000000111110,  // 0.4862793982028961
14'b00000000101111,  // 0.37162142992019653
14'b00000000111010,  // 0.45989668369293213
14'b00000010100110,  // 1.2998151779174805
14'b11111101111101,  // -1.016528844833374
14'b11111111010010,  // -0.35249894857406616
14'b00000000111001,  // 0.44582197070121765
14'b11111111110001,  // -0.1119980737566948
14'b11111111110111,  // -0.06717441976070404
14'b00000000000000,  // 0.00487547367811203
14'b00000000011000,  // 0.1946917623281479
14'b11111110011100,  // -0.7796769738197327
14'b00000001011101,  // 0.7287401556968689
14'b00000011011011,  // 1.714877724647522
14'b11111100110011,  // -1.5971007347106934
14'b00000000001001,  // 0.07393483817577362
14'b00000000101001,  // 0.3225609362125397
14'b00000001101100,  // 0.8453295230865479
14'b00000001110011,  // 0.898597240447998
14'b00000000100000,  // 0.2548799514770508
14'b00000001111100,  // 0.9735668301582336
14'b00000010010000,  // 1.1261906623840332
14'b00000000111001,  // 0.44768181443214417
14'b11111011010000   // -2.3676068782806396
};
endpackage