// Width: 24
// NFRAC: 12
package dense_4_24_12;

localparam logic signed [23:0] weights [32][5] = '{ 
{24'b111111111111111111001111, 24'b000000000000010100001100, 24'b111111111111101100111011, 24'b000000000000000100001101, 24'b111111111111111001001100}, 
{24'b111111111111011100010011, 24'b111111111111111100011110, 24'b000000000000011101011101, 24'b111111111111111111001101, 24'b000000000000000001000100}, 
{24'b000000000000010111110001, 24'b000000000000001101100011, 24'b111111111111111110001101, 24'b111111111111100110000011, 24'b111111111111110010100000}, 
{24'b111111111111100111111101, 24'b111111111111101000001000, 24'b111111111111111000110110, 24'b000000000000010011101100, 24'b000000000000001111000010}, 
{24'b000000000000000111110100, 24'b000000000000001000001111, 24'b000000000000001010000011, 24'b111111111111111110110101, 24'b111111111110111111001011}, 
{24'b000000000000010100111011, 24'b111111111111100110110000, 24'b000000000000001011100111, 24'b111111111111110101101011, 24'b111111111111110101000110}, 
{24'b111111111111100110010100, 24'b000000000000000010010001, 24'b111111111111111111111111, 24'b000000000000001011001001, 24'b000000000000000100011010}, 
{24'b111111111111111111111000, 24'b000000000000010010001101, 24'b111111111111100110111010, 24'b000000000000001010011010, 24'b000000000000001000101101}, 
{24'b000000000000001010011101, 24'b111111111111110101001010, 24'b000000000000000000000101, 24'b111111111111100010011101, 24'b111111111111110000000101}, 
{24'b111111111111111111111111, 24'b111111111111101110111101, 24'b000000000000001011011000, 24'b000000000000011011100001, 24'b000000000000000000000000}, 
{24'b111111111111110111101011, 24'b111111111111110110101111, 24'b000000000000000000000000, 24'b000000000000100101001101, 24'b111111111111101110110111}, 
{24'b000000000000001010110101, 24'b000000000000001110101010, 24'b111111111111101010001111, 24'b111111111111111110001111, 24'b000000000000000111110010}, 
{24'b000000000000000000000000, 24'b000000000000001010101110, 24'b000000000000000000100100, 24'b111111111111110010101100, 24'b111111111111011000001000}, 
{24'b000000000000001011010110, 24'b000000000000000100000101, 24'b000000000000011010110110, 24'b111111111111111011100001, 24'b111111111111100100100111}, 
{24'b000000000000000101110011, 24'b111111111111111100111010, 24'b111111111111101000111011, 24'b111111111111111101111000, 24'b000000000000100010010100}, 
{24'b111111111111100001101010, 24'b111111111111110000010111, 24'b111111111111110001110000, 24'b000000000000011001100001, 24'b000000000000000010000011}, 
{24'b000000000000010110001000, 24'b111111111111110101000000, 24'b111111111111110111010100, 24'b111111111111110001100011, 24'b111111111111111100001010}, 
{24'b000000000000001100011110, 24'b111111111111111101011010, 24'b111111111111100101100111, 24'b111111111111111110000010, 24'b000000000000000100100001}, 
{24'b000000000000010000100010, 24'b000000000000000010101010, 24'b111111111111110010000011, 24'b000000000000000000000000, 24'b111111111111100111111100}, 
{24'b000000000000001110110011, 24'b111111111111111010011101, 24'b111111111111110010011000, 24'b000000000000001101010000, 24'b000000000000000110000101}, 
{24'b000000000000000100010101, 24'b111111111111111110000011, 24'b000000000000010011000010, 24'b111111111111100100011010, 24'b111111111111111110101000}, 
{24'b000000000000000000000000, 24'b000000000000000111100010, 24'b000000000000011111001001, 24'b111111111111011110110101, 24'b111111111111011000011110}, 
{24'b111111111111111001101101, 24'b000000000000000111000001, 24'b000000000000001011010101, 24'b111111111111101001001010, 24'b000000000000100001011011}, 
{24'b111111111111111111111110, 24'b000000000000001010100011, 24'b000000000000010010000101, 24'b000000000000000010011011, 24'b111111111111011011011000}, 
{24'b111111111111110101001010, 24'b000000000000010111010100, 24'b111111111111110001101100, 24'b000000000000000000010111, 24'b000000000000011000110101}, 
{24'b000000000000000001101011, 24'b000000000000010001000000, 24'b000000000000000001111001, 24'b111111111111010000001000, 24'b000000000000100011000101}, 
{24'b111111111111100010100101, 24'b111111111111110000011010, 24'b000000000000001101101101, 24'b000000000000001111101001, 24'b000000000000001100111010}, 
{24'b000000000000000000010000, 24'b000000000000001111011011, 24'b111111111111111101101010, 24'b111111111111110110010111, 24'b000000000000000010000001}, 
{24'b111111111111111001010101, 24'b000000000000001111110000, 24'b111111111111011111110000, 24'b000000000000001000111000, 24'b111111111111110101110111}, 
{24'b111111111111111110110100, 24'b000000000000001001000010, 24'b111111111111110101001100, 24'b111111111111100110010111, 24'b000000000000100101111111}, 
{24'b000000000000011100101110, 24'b000000000000000100011110, 24'b000000000000010100110001, 24'b111111111111011010010000, 24'b111111111111101011110101}, 
{24'b111111111111111100001101, 24'b111111111111100111010010, 24'b000000000000010111011010, 24'b000000000000000100100010, 24'b000000000000001000001010}
};

localparam logic signed [23:0] bias [5] = '{
24'b111111111111111100000001,  // -0.06223141402006149
24'b111111111111111011111111,  // -0.06270556896924973
24'b111111111111111011100000,  // -0.07014333456754684
24'b000000000000000101010000,  // 0.0820775106549263
24'b000000000000001101110010   // 0.2155742198228836
};
endpackage