// Width: 25
// NFRAC: 12
package dense_3_25_13;

localparam logic signed [24:0] weights [32][32] = '{ 
{25'b1111111111111111100110110, 25'b1111111111111100100000001, 25'b1111111111111100110000010, 25'b1111111111111110011110011, 25'b0000000000000010101111101, 25'b0000000000000000010110011, 25'b1111111111111111111001011, 25'b1111111111111111111111100, 25'b1111111111111111111111111, 25'b1111111111111111111111111, 25'b0000000000000001000000100, 25'b1111111111111011110010001, 25'b1111111111111111100001011, 25'b0000000000000110110001101, 25'b1111111111111110000100010, 25'b1111111111111000100010011, 25'b1111111111111111101101011, 25'b0000000000000000111001000, 25'b0000000000000011011110101, 25'b1111111111111101001101101, 25'b1111111111110111011110011, 25'b1111111111111111101000011, 25'b0000000000000000011001001, 25'b1111111111111100110001100, 25'b0000000000000000000000000, 25'b0000000000001000000110011, 25'b1111111111110100010110010, 25'b1111111111111110001110100, 25'b1111111111111100111001000, 25'b1111111111111110110011001, 25'b0000000000000011011000100, 25'b1111111111111110101110011}, 
{25'b0000000000000101111110110, 25'b0000000000001101110101110, 25'b0000000000000011001101110, 25'b1111111111111010101111010, 25'b0000000000000001111101000, 25'b1111111111111101110100000, 25'b1111111111111111001000011, 25'b0000000000001000101110000, 25'b0000000000000000000011000, 25'b1111111111111111111111111, 25'b1111111111111111101111101, 25'b1111111111111011010010110, 25'b1111111111111110011000111, 25'b0000000000000100010100101, 25'b1111111111101111001001110, 25'b1111111111111100001110101, 25'b1111111111111111111111111, 25'b1111111111111111111011110, 25'b1111111111111111100101000, 25'b1111111111111110101011111, 25'b1111111111111101111011101, 25'b1111111111111101110011000, 25'b0000000000000000001000110, 25'b1111111111111111111111001, 25'b1111111111111111111100101, 25'b1111111111110111011011000, 25'b0000000000000000000110000, 25'b0000000000000011110001001, 25'b1111111111111111011111100, 25'b1111111111111010011110110, 25'b0000000000000000000001011, 25'b0000000000000000010011011}, 
{25'b1111111111111000000111100, 25'b0000000000000001011110010, 25'b0000000000000000000101011, 25'b0000000000000010100101001, 25'b1111111111111010111101010, 25'b0000000000000000000000010, 25'b0000000000000000000000110, 25'b1111111111111001010010010, 25'b0000000000000100010010011, 25'b1111111111111101111001110, 25'b1111111111111101111011001, 25'b1111111111110100000110101, 25'b1111111111111101100000110, 25'b0000000000000100000101100, 25'b0000000000000010000111000, 25'b1111111111111111111111001, 25'b1111111111111111000101011, 25'b1111111111111111110011111, 25'b1111111111111001011110111, 25'b0000000000000000000001100, 25'b0000000000000000111111110, 25'b0000000000000000100011010, 25'b0000000000000001101011000, 25'b0000000000000111000010100, 25'b0000000000000000010011011, 25'b1111111111111001101100011, 25'b0000000000000110001000111, 25'b0000000000000000000000010, 25'b0000000000000001010100111, 25'b1111111111111111110100101, 25'b0000000000000000000000011, 25'b0000000000010010001001101}, 
{25'b0000000000000110101100111, 25'b1111111111111111111111111, 25'b1111111111111110011100011, 25'b0000000000001010011110000, 25'b0000000000001001110100110, 25'b0000000000000000000000001, 25'b0000000000000000100101101, 25'b0000000000000110100000101, 25'b1111111111111100110101010, 25'b1111111111111111111111111, 25'b1111111111111001011010011, 25'b0000000000000000111101010, 25'b0000000000000010001000011, 25'b1111111111111010000001010, 25'b0000000000000000101111111, 25'b1111111111111110101110001, 25'b1111111111111111111111111, 25'b1111111111111101000101100, 25'b0000000000000000010011101, 25'b0000000000000000011100010, 25'b0000000000000000001000001, 25'b1111111111111111011010101, 25'b0000000000001001100011001, 25'b0000000000000101011111000, 25'b0000000000000101010001010, 25'b0000000000000011111110001, 25'b0000000000000101011101110, 25'b0000000000000000000000001, 25'b1111111111111111000011100, 25'b0000000000000111001111111, 25'b0000000000000011111111100, 25'b1111111111111110100110000}, 
{25'b0000000000001000000000010, 25'b1111111111111111010000001, 25'b1111111111111010011101000, 25'b1111111111110011111110011, 25'b0000000000000111101000111, 25'b0000000000000000000000001, 25'b1111111111111001011011111, 25'b1111111111111011011110100, 25'b1111111111111111010000010, 25'b1111111111110011000011010, 25'b1111111111101110010100101, 25'b0000000000000111100100000, 25'b0000000000001010101100110, 25'b0000000000001000010111111, 25'b1111111111110110110011001, 25'b1111111111110011100110011, 25'b0000000000000000000000000, 25'b1111111111111101101111001, 25'b0000000000000011001101100, 25'b0000000000000010001110000, 25'b1111111111111100111111000, 25'b1111111111111111111001011, 25'b0000000000001011100010111, 25'b1111111111101010000000010, 25'b0000000000000001011010001, 25'b1111111111110101011101101, 25'b0000000000000001000011000, 25'b1111111111111100000001111, 25'b1111111111111011001110011, 25'b1111111111111111111111101, 25'b0000000000000001000111101, 25'b0000000000001001010010011}, 
{25'b0000000000000000101100001, 25'b1111111111111111010101101, 25'b1111111111111011000101100, 25'b1111111111111011110101011, 25'b0000000000000101111100101, 25'b0000000000000000000000001, 25'b1111111111111011100001100, 25'b1111111111111101110100100, 25'b1111111111111001001001100, 25'b1111111111111110111110011, 25'b1111111111111111111111100, 25'b0000000000000010100100001, 25'b0000000000000000000000000, 25'b0000000000000101101110010, 25'b1111111111110111111010000, 25'b1111111111111101111101010, 25'b0000000000000001011011001, 25'b1111111111111011010011111, 25'b1111111111111100110101101, 25'b1111111111111111111111111, 25'b0000000000000000001100011, 25'b0000000000000100110010110, 25'b0000000000000111011110001, 25'b1111111111111111110101000, 25'b1111111111111111111111100, 25'b0000000000000110011010010, 25'b1111111111110111001101010, 25'b1111111111111111111111111, 25'b1111111111111100001101110, 25'b1111111111111111011010010, 25'b1111111111111111111100110, 25'b0000000000000000000110101}, 
{25'b0000000000000001000010101, 25'b1111111111111010101011100, 25'b0000000000000001101110111, 25'b1111111111111111011000100, 25'b1111111111111111111000010, 25'b0000000000000010011011000, 25'b1111111111111110010011011, 25'b1111111111110101001010101, 25'b1111111111111111111111111, 25'b1111111111111100101010101, 25'b1111111111111000101100010, 25'b0000000000000111100011100, 25'b0000000000000000000111010, 25'b0000000000001010111100110, 25'b0000000000001101010000100, 25'b0000000000000000000010101, 25'b1111111111111111111111111, 25'b1111111111111010111101001, 25'b1111111111111111000000100, 25'b0000000000000100010111111, 25'b1111111111110011111111111, 25'b0000000000000010011111101, 25'b0000000000000101001110001, 25'b0000000000000000010011011, 25'b0000000000000010011001101, 25'b0000000000010011111001001, 25'b1111111111111001101100011, 25'b1111111111111110100011001, 25'b1111111111111100111101100, 25'b0000000000000111110010110, 25'b1111111111111111001101101, 25'b1111111111111101010010100}, 
{25'b1111111111110110011101011, 25'b0000000000000000011000011, 25'b1111111111110101111011101, 25'b0000000000000110111101101, 25'b0000000000010000011100101, 25'b0000000000000001110110111, 25'b0000000000000000000011111, 25'b0000000000000000110000010, 25'b1111111111111111111111111, 25'b0000000000000010000011000, 25'b0000000000010100110100010, 25'b1111111111111111111111101, 25'b0000000000000110000110010, 25'b0000000000001001111101111, 25'b0000000000001100010011000, 25'b0000000000010000110011010, 25'b0000000000000000000000000, 25'b1111111111111000010110011, 25'b0000000000000101011000010, 25'b1111111111111111111010011, 25'b1111111111110101110010110, 25'b1111111111111100010111101, 25'b0000000000000000001101110, 25'b1111111111111110101011001, 25'b1111111111110111111110101, 25'b0000000000011110000000100, 25'b1111111111111100011111001, 25'b0000000000000000000000000, 25'b0000000000000000000000000, 25'b0000000000001110001000001, 25'b0000000000000001011010110, 25'b0000000000000110010001001}, 
{25'b0000000000000110110000011, 25'b1111111111111111101100000, 25'b0000000000000000000000010, 25'b1111111111111111010011101, 25'b0000000000000001010011100, 25'b1111111111111111011001000, 25'b1111111111111111111111101, 25'b0000000000000010100000101, 25'b0000000000000011011000011, 25'b1111111111111011100111011, 25'b0000000000000010001111011, 25'b0000000000000010111111111, 25'b0000000000000000001100001, 25'b0000000000000101010100110, 25'b1111111111111100011001100, 25'b1111111111110011001111111, 25'b0000000000000000000000000, 25'b1111111111111111110001101, 25'b1111111111111111100100101, 25'b1111111111111000000001011, 25'b1111111111111111111110110, 25'b0000000000000000000000000, 25'b1111111111111100110000011, 25'b1111111111111111110001100, 25'b1111111111111110011110101, 25'b0000000000000010011111100, 25'b0000000000000101111110101, 25'b1111111111111110000101101, 25'b1111111111111111001101101, 25'b1111111111111111010110110, 25'b0000000000000000011011101, 25'b1111111111111001101110001}, 
{25'b1111111111111101001010000, 25'b0000000000000110001001101, 25'b0000000000000000000000000, 25'b0000000000000000000000000, 25'b0000000000001100101011010, 25'b0000000000000101001001111, 25'b1111111111111111111111111, 25'b1111111111110111000111100, 25'b0000000000000001111000101, 25'b1111111111110100110101101, 25'b1111111111101001100011001, 25'b1111111111111111111111111, 25'b0000000000000000000000010, 25'b0000000000000110110111010, 25'b0000000000000001110001101, 25'b0000000000000000000000000, 25'b1111111111111010101111101, 25'b0000000000000000000000010, 25'b0000000000000000000110111, 25'b0000000000000000111110000, 25'b0000000000000011111001101, 25'b1111111111111111100101111, 25'b1111111111111010001111001, 25'b0000000000000000001000011, 25'b1111111111111111110100011, 25'b0000000000010001010011011, 25'b0000000000000101001110011, 25'b1111111111111111111111100, 25'b1111111111111110110111011, 25'b0000000000001010101100010, 25'b1111111111111111010111001, 25'b1111111111111110100110010}, 
{25'b1111111111110111101000011, 25'b0000000000000010110011011, 25'b1111111111111111011100011, 25'b1111111111111111111111111, 25'b1111111111111100000011111, 25'b1111111111111001111101010, 25'b0000000000000000110001001, 25'b0000000000000010010011101, 25'b1111111111111111111111111, 25'b1111111111111101010000101, 25'b1111111111110110110101101, 25'b0000000000000011001101101, 25'b0000000000000100110111011, 25'b0000000000000000000000000, 25'b0000000000001101011011000, 25'b1111111111110111000000110, 25'b0000000000000001101010011, 25'b1111111111111001101111100, 25'b0000000000000100100000110, 25'b1111111111111111111111110, 25'b1111111111111111011000100, 25'b0000000000000001000111111, 25'b0000000000000001111101101, 25'b0000000000000000000000001, 25'b1111111111111000000110011, 25'b0000000000000000011111110, 25'b1111111111110111000011110, 25'b1111111111111111010111010, 25'b1111111111111111111111110, 25'b0000000000001010110011111, 25'b1111111111111100111101010, 25'b0000000000000000000000010}, 
{25'b1111111111111111111111111, 25'b0000000000000001110101100, 25'b0000000000000000000000010, 25'b0000000000000110010000101, 25'b1111111111111110001000000, 25'b1111111111111111010011111, 25'b0000000000000000111011111, 25'b1111111111111111111010000, 25'b1111111111111111010000100, 25'b0000000000001010010000000, 25'b0000000000001011001011111, 25'b0000000000000000000000101, 25'b1111111111111010101011011, 25'b1111111111110100110000111, 25'b1111111111111111001100000, 25'b0000000000000000000000001, 25'b0000000000000000000000001, 25'b1111111111111110111110110, 25'b1111111111111000011000000, 25'b0000000000000110000111100, 25'b0000000000000000000010001, 25'b0000000000000101111011111, 25'b1111111111111111111111110, 25'b0000000000001000111111111, 25'b0000000000000001111110101, 25'b0000000000000100111001101, 25'b0000000000000111010010011, 25'b1111111111111111001011000, 25'b1111111111111001101111001, 25'b1111111111111000111100110, 25'b1111111111111111111010110, 25'b1111111111110101010011000}, 
{25'b1111111111111100011000001, 25'b1111111111111111111111111, 25'b0000000000000001111010001, 25'b1111111111111001010011000, 25'b0000000000000001011000001, 25'b1111111111111111111111111, 25'b1111111111111100100001100, 25'b1111111111111111110110001, 25'b1111111111111101111111100, 25'b0000000000000000100110000, 25'b0000000000000001001111110, 25'b1111111111111110110110110, 25'b0000000000000000010000111, 25'b0000000000000011000000001, 25'b1111111111110101111111111, 25'b1111111111111100000101011, 25'b0000000000000011101001101, 25'b1111111111111101001010110, 25'b0000000000000000000000000, 25'b1111111111111111100110010, 25'b0000000000000011000101100, 25'b0000000000000000001000001, 25'b1111111111111111100000001, 25'b0000000000000000101011100, 25'b0000000000000100010011111, 25'b1111111111111110010101100, 25'b0000000000000000000000001, 25'b1111111111111000110001011, 25'b1111111111111100110111100, 25'b1111111111111111111000110, 25'b0000000000000010110001100, 25'b0000000000000000000000010}, 
{25'b1111111111110111101011110, 25'b0000000000000110101110011, 25'b1111111111111111111111111, 25'b1111111111111111111001001, 25'b1111111111111111110110001, 25'b0000000000000010110011100, 25'b1111111111111111111111110, 25'b0000000000001100010110100, 25'b1111111111111111110000110, 25'b1111111111111111111111111, 25'b0000000000000011010010110, 25'b0000000000000000101001111, 25'b0000000000000000000110101, 25'b0000000000000000000000001, 25'b0000000000000001111100101, 25'b0000000000000101010010000, 25'b0000000000000010110110011, 25'b0000000000000010101010101, 25'b1111111111111111110111010, 25'b0000000000000100111010100, 25'b0000000000000001100111000, 25'b0000000000000000101001011, 25'b1111111111111111110111001, 25'b0000000000000100000100000, 25'b1111111111111110011010000, 25'b1111111111111010100100111, 25'b1111111111111110100001011, 25'b1111111111111111111111111, 25'b0000000000000001101000000, 25'b0000000000000000011110011, 25'b0000000000000011001000000, 25'b0000000000000111101010101}, 
{25'b1111111111111111101100111, 25'b1111111111111001110001010, 25'b0000000000000000110100111, 25'b1111111111111111111111000, 25'b0000000000001110101010000, 25'b1111111111111100101011101, 25'b1111111111110110110110101, 25'b0000000000000000000000001, 25'b0000000000000000000000000, 25'b1111111111111111100101100, 25'b0000000000000000110001100, 25'b0000000000000110111111001, 25'b0000000000000101001001101, 25'b0000000000000000001010111, 25'b0000000000000000100010001, 25'b1111111111111101001101000, 25'b0000000000000000100010001, 25'b1111111111111111011001001, 25'b0000000000000000000000000, 25'b0000000000000001001101001, 25'b1111111111111111011001101, 25'b0000000000000000010011100, 25'b0000000000000100010000101, 25'b0000000000000000100101110, 25'b1111111111111111110011101, 25'b1111111111111001011001011, 25'b0000000000000011010000000, 25'b1111111111111111111111111, 25'b1111111111111111111111101, 25'b1111111111111110010011001, 25'b1111111111111111101010000, 25'b1111111111111110111111111}, 
{25'b0000000000000000000111010, 25'b1111111111111110111111001, 25'b1111111111111101111110111, 25'b1111111111111100100000000, 25'b1111111111110111010000010, 25'b0000000000001001110000000, 25'b0000000000000000000000001, 25'b0000000000000010101100111, 25'b0000000000000100100101111, 25'b0000000000000000001101001, 25'b1111111111111111011101010, 25'b0000000000000111100111000, 25'b0000000000000011100101001, 25'b1111111111111010001001101, 25'b1111111111111101011001110, 25'b1111111111111111010101110, 25'b1111111111111001101000000, 25'b1111111111111111101110001, 25'b0000000000000000000000001, 25'b1111111111111111111011010, 25'b0000000000000010011111101, 25'b1111111111111101110011111, 25'b0000000000000000000000000, 25'b0000000000000001001110110, 25'b1111111111111111111111111, 25'b1111111111111010100010000, 25'b0000000000000010100000011, 25'b0000000000000000000000011, 25'b0000000000000000101101101, 25'b0000000000000000001011001, 25'b1111111111111010111100010, 25'b0000000000000000010101010}, 
{25'b1111111111111100110111001, 25'b1111111111111101011110110, 25'b0000000000000001001110010, 25'b1111111111111110000000111, 25'b1111111111111110100100000, 25'b0000000000000001110110111, 25'b1111111111111111111010110, 25'b0000000000000000100011110, 25'b0000000000000010000110001, 25'b1111111111111111111111101, 25'b0000000000000001111110101, 25'b1111111111111101111101101, 25'b1111111111111111110110000, 25'b1111111111111111111111110, 25'b0000000000000001101001111, 25'b1111111111111111111111111, 25'b0000000000000111110100001, 25'b1111111111111111101110001, 25'b0000000000000011111110000, 25'b1111111111111101010010001, 25'b0000000000000010100010000, 25'b0000000000000001000000010, 25'b0000000000000001010110011, 25'b0000000000000000100101001, 25'b1111111111111110101100101, 25'b1111111111111011100010100, 25'b1111111111111011110110101, 25'b0000000000000001101110100, 25'b1111111111111110101010010, 25'b0000000000000000000000100, 25'b1111111111111111100011111, 25'b0000000000000011101101101}, 
{25'b1111111111111111111111111, 25'b1111111111111001100001011, 25'b1111111111111001101001111, 25'b1111111111111111111111111, 25'b0000000000001010000110011, 25'b1111111111111110100011000, 25'b0000000000000000000000001, 25'b0000000000000111101110111, 25'b1111111111111101101000111, 25'b0000000000000000000000000, 25'b1111111111111001010100010, 25'b1111111111111000001010000, 25'b0000000000000111001011000, 25'b0000000000000010011010110, 25'b1111111111111110000011110, 25'b1111111111111011100111101, 25'b0000000000000010110000100, 25'b0000000000000000000000011, 25'b1111111111111100001100100, 25'b0000000000000000011011001, 25'b0000000000000001000111001, 25'b1111111111111110100101011, 25'b0000000000000100100010110, 25'b1111111111110000010100110, 25'b0000000000000000101001111, 25'b0000000000000011110100110, 25'b1111111111111111010101110, 25'b0000000000000000001111010, 25'b1111111111111100010001001, 25'b1111111111111111111111110, 25'b1111111111111100110010000, 25'b1111111111111111100111010}, 
{25'b0000000000000011011001101, 25'b0000000000000101100001011, 25'b0000000000001000110011111, 25'b1111111111111100101110100, 25'b0000000000000110101010000, 25'b0000000000000100111001101, 25'b0000000000000000000000100, 25'b0000000000000111010010011, 25'b0000000000000101101101101, 25'b1111111111111110010010100, 25'b0000000000001011001110011, 25'b1111111111111010011010011, 25'b0000000000001001111100010, 25'b0000000000000111001001000, 25'b1111111111101110110101010, 25'b1111111111111111111111000, 25'b0000000000000000000000000, 25'b0000000000000000000101111, 25'b0000000000000100001010001, 25'b1111111111110111111100101, 25'b0000000000000011100010111, 25'b1111111111111100100110111, 25'b1111111111111000001001111, 25'b1111111111111101011111011, 25'b0000000000000101010001010, 25'b1111111111110101011100011, 25'b1111111111111010101110010, 25'b1111111111111111010101110, 25'b1111111111111111111111110, 25'b1111111111110110111110001, 25'b0000000000000110010100111, 25'b0000000000000000000000011}, 
{25'b1111111111111111001101100, 25'b0000000000000000000000101, 25'b1111111111111111111111111, 25'b1111111111111111111111111, 25'b1111111111111010011000011, 25'b0000000000000000001001011, 25'b0000000000000000001000011, 25'b1111111111111111110000100, 25'b1111111111111111100111001, 25'b1111111111111111010000111, 25'b0000000000000010001110010, 25'b1111111111111111111111001, 25'b0000000000000001010100111, 25'b1111111111111010100001100, 25'b0000000000000001101101011, 25'b1111111111111111111111010, 25'b0000000000000010010000000, 25'b0000000000000111001010011, 25'b1111111111111010010110110, 25'b0000000000000000110101001, 25'b1111111111111110011010100, 25'b0000000000000010000011101, 25'b0000000000000011000010101, 25'b1111111111111110101000101, 25'b1111111111111011111110110, 25'b0000000000000000010101000, 25'b0000000000001101010001001, 25'b1111111111111111100111001, 25'b1111111111111111110000010, 25'b0000000000000101001100000, 25'b0000000000000000000000001, 25'b0000000000001101110010101}, 
{25'b1111111111110111101001111, 25'b0000000000000000100101000, 25'b1111111111111100100010011, 25'b0000000000000110001000000, 25'b0000000000000001110000010, 25'b1111111111111111011111101, 25'b1111111111111111111111111, 25'b1111111111111111111111111, 25'b1111111111111011001001100, 25'b1111111111111111011110001, 25'b0000000000000000000000001, 25'b1111111111110111000111011, 25'b0000000000000000001100110, 25'b1111111111111111010111010, 25'b1111111111111111111101011, 25'b1111111111111111111111110, 25'b1111111111111110001000100, 25'b0000000000000000000101100, 25'b0000000000000000000011001, 25'b0000000000000010100010011, 25'b0000000000000000010001111, 25'b0000000000000000000000000, 25'b0000000000000000000000001, 25'b1111111111111111110111101, 25'b0000000000000000000000010, 25'b0000000000000000010010110, 25'b0000000000001001010011010, 25'b1111111111111111111111111, 25'b1111111111111111111111110, 25'b1111111111111111010110010, 25'b0000000000000010110011010, 25'b1111111111111111100101111}, 
{25'b1111111111111111111110011, 25'b1111111111111101100101000, 25'b0000000000000011010001001, 25'b0000000000000000101000111, 25'b1111111111111010000011010, 25'b0000000000000000000000100, 25'b0000000000000100100100110, 25'b1111111111111111111111110, 25'b0000000000000000000000000, 25'b1111111111111110011011000, 25'b0000000000000001110101101, 25'b0000000000000000010011011, 25'b0000000000000101001011010, 25'b1111111111110111001110100, 25'b1111111111111110011111001, 25'b1111111111111111101110011, 25'b0000000000000011011101010, 25'b1111111111111001110110101, 25'b0000000000000000010101110, 25'b1111111111110011111011010, 25'b1111111111111111101100101, 25'b1111111111111110000110001, 25'b1111111111111111010110101, 25'b0000000000000100101110110, 25'b1111111111111110110011101, 25'b1111111111111011100000001, 25'b0000000000000001011100100, 25'b0000000000000000000000010, 25'b0000000000000110010101010, 25'b0000000000001000010111110, 25'b1111111111111010110000000, 25'b1111111111111000110100000}, 
{25'b0000000000000001000101000, 25'b0000000000000000011010001, 25'b1111111111111001010111111, 25'b1111111111111111000101111, 25'b1111111111111111111111111, 25'b0000000000000000000010001, 25'b0000000000000001101100110, 25'b0000000000000110100101001, 25'b0000000000000000000000000, 25'b0000000000000000010100110, 25'b0000000000000001000111101, 25'b1111111111110111010111101, 25'b1111111111111110111011110, 25'b1111111111110110010101110, 25'b0000000000000111101100011, 25'b0000000000000000000000011, 25'b1111111111111111111111001, 25'b1111111111110101101111110, 25'b1111111111111111111111101, 25'b1111111111111110110011110, 25'b1111111111111111101010101, 25'b0000000000000000000000000, 25'b0000000000000000111111110, 25'b1111111111111101100110000, 25'b0000000000000000110110011, 25'b0000000000000110100100110, 25'b0000000000000110110100101, 25'b0000000000000110001111111, 25'b0000000000000100111011011, 25'b0000000000000000000000001, 25'b0000000000000001110100111, 25'b0000000000001100100010010}, 
{25'b1111111111111111100110001, 25'b1111111111111100001100011, 25'b0000000000000110001110101, 25'b1111111111111110010110101, 25'b0000000000000001000111011, 25'b0000000000000010101011111, 25'b1111111111111111111111111, 25'b1111111111111011011010001, 25'b1111111111111110101000110, 25'b1111111111110110011000110, 25'b0000000000000111001010000, 25'b0000000000000000000011111, 25'b0000000000000110101101001, 25'b0000000000001010101110001, 25'b1111111111111110001000110, 25'b1111111111110010000100011, 25'b1111111111111110010101101, 25'b0000000000000111100001001, 25'b1111111111111011011110010, 25'b1111111111111100101010010, 25'b0000000000000000111100110, 25'b0000000000000000000001000, 25'b1111111111110111010001111, 25'b1111111111111100111100001, 25'b1111111111111111010111110, 25'b1111111111111110000011010, 25'b0000000000000001110010111, 25'b0000000000001011010000011, 25'b0000000000000011111011011, 25'b1111111111111111111111111, 25'b0000000000000001010010101, 25'b0000000000000000011100010}, 
{25'b0000000000000000101011011, 25'b0000000000000111010000100, 25'b0000000000000000000000000, 25'b0000000000000100101110100, 25'b0000000000001101010011001, 25'b1111111111111101010001001, 25'b1111111111111111111111111, 25'b1111111111111111010010101, 25'b0000000000000100101100000, 25'b1111111111111100111011111, 25'b1111111111111111111110101, 25'b0000000000000101010101010, 25'b0000000000000000001000101, 25'b0000000000000000011100000, 25'b1111111111100111100100010, 25'b1111111111111110101110101, 25'b0000000000000000000000000, 25'b0000000000000011001101100, 25'b1111111111111111111100100, 25'b0000000000000100110001110, 25'b1111111111111111111111110, 25'b1111111111111101001111000, 25'b1111111111110111000000100, 25'b0000000000000010000101111, 25'b0000000000000100100100110, 25'b1111111111101110010000001, 25'b1111111111111111111111110, 25'b0000000000000000000000001, 25'b0000000000001000101101001, 25'b1111111111110011001011011, 25'b0000000000000000000001110, 25'b1111111111111111111001110}, 
{25'b0000000000000000001001101, 25'b1111111111111010100100001, 25'b0000000000000000110111010, 25'b1111111111111111110000101, 25'b0000000000000000110101010, 25'b0000000000001000011101110, 25'b1111111111110100011001110, 25'b0000000000000000100011001, 25'b0000000000000110110001100, 25'b1111111111111010100110101, 25'b1111111111111111101000001, 25'b0000000000000000110010000, 25'b1111111111111111110110110, 25'b0000000000000010110111001, 25'b0000000000000001101101111, 25'b1111111111111111101110111, 25'b0000000000000001000100101, 25'b0000000000000000000000010, 25'b0000000000000000010110000, 25'b0000000000000110000100111, 25'b1111111111111111100011010, 25'b1111111111111000010000000, 25'b1111111111110110010100100, 25'b1111111111111100111001101, 25'b1111111111110110100011001, 25'b0000000000000011010101000, 25'b0000000000001001111110001, 25'b0000000000000101111001100, 25'b1111111111111111110101010, 25'b1111111111111010000010011, 25'b1111111111111011000001110, 25'b0000000000000000111101001}, 
{25'b0000000000000000110101001, 25'b1111111111111000010110111, 25'b1111111111111111101110101, 25'b0000000000000010011010000, 25'b1111111111111000010110000, 25'b0000000000000010101101110, 25'b1111111111111111111111111, 25'b1111111111111111111111110, 25'b1111111111111111111111111, 25'b0000000000000000000000001, 25'b0000000000000100001110101, 25'b1111111111111111101110010, 25'b0000000000000000001001111, 25'b0000000000000000000000010, 25'b0000000000000010000010011, 25'b1111111111111111101110101, 25'b0000000000000000000010110, 25'b1111111111111111111111010, 25'b1111111111111010110110001, 25'b1111111111110111111010001, 25'b1111111111111111111111011, 25'b1111111111110111011101010, 25'b1111111111111011001011100, 25'b1111111111111010000011010, 25'b0000000000001110001111111, 25'b0000000000000000010010000, 25'b1111111111111111010000110, 25'b0000000000000101000100111, 25'b0000000000001110010111000, 25'b0000000000000110010100010, 25'b1111111111101111000010000, 25'b1111111111111101000010000}, 
{25'b0000000000000110000000111, 25'b1111111111111111111111100, 25'b0000000000000100000001000, 25'b1111111111111111101011101, 25'b0000000000000111101111010, 25'b1111111111111101101101111, 25'b0000000000000001001000100, 25'b0000000000000110101100010, 25'b0000000000000100010010001, 25'b1111111111110111101001010, 25'b1111111111111111000000111, 25'b0000000000000001111101110, 25'b0000000000000001000110100, 25'b1111111111111111110001000, 25'b0000000000000001010110111, 25'b0000000000000000000000010, 25'b0000000000000101110011000, 25'b0000000000000000100011111, 25'b0000000000000101111111001, 25'b1111111111111110111100111, 25'b1111111111111101111101100, 25'b1111111111111110110011011, 25'b1111111111111111111111110, 25'b0000000000000100110101000, 25'b1111111111111100110000110, 25'b1111111111111111111001101, 25'b0000000000000000000000000, 25'b0000000000000000000000010, 25'b0000000000000000000000001, 25'b0000000000000100101011000, 25'b1111111111111010110111101, 25'b1111111111111111101000001}, 
{25'b1111111111111111111111010, 25'b1111111111111111100000011, 25'b1111111111111000100011110, 25'b0000000000000100100011010, 25'b0000000000000011100100100, 25'b1111111111111110001111110, 25'b1111111111111111111111110, 25'b1111111111111100010111101, 25'b0000000000000000000110111, 25'b1111111111111111111111101, 25'b1111111111111011001011011, 25'b1111111111111100000011110, 25'b0000000000000111101010100, 25'b0000000000000000000000000, 25'b1111111111111101111101001, 25'b1111111111111111111111111, 25'b0000000000000011011011001, 25'b1111111111111111111111110, 25'b1111111111111111111111111, 25'b1111111111111100100010110, 25'b0000000000000101000011111, 25'b0000000000000000000000000, 25'b0000000000000010011111111, 25'b1111111111111111100010101, 25'b0000000000000010100000110, 25'b0000000000000000000010010, 25'b0000000000000000000000000, 25'b0000000000000011110110100, 25'b1111111111111100111011010, 25'b1111111111111111010000110, 25'b0000000000000010100100011, 25'b1111111111111110010011100}, 
{25'b1111111111111111101110110, 25'b1111111111111011000100000, 25'b0000000000001001100000101, 25'b1111111111111110111101011, 25'b0000000000000011001001000, 25'b1111111111111011011011000, 25'b0000000000000000000000000, 25'b0000000000000000100011000, 25'b1111111111111000010101011, 25'b1111111111111111110010111, 25'b1111111111111110000001010, 25'b0000000000000000111011100, 25'b1111111111111010110000001, 25'b0000000000000010001101001, 25'b0000000000000011001111001, 25'b0000000000000001110000001, 25'b0000000000000001010111110, 25'b1111111111111111011001000, 25'b1111111111110100101010110, 25'b1111111111111111110010001, 25'b1111111111111111000101101, 25'b0000000000000010001111001, 25'b1111111111111110001110010, 25'b1111111111111111111111111, 25'b0000000000000011001010011, 25'b1111111111111111010001010, 25'b1111111111111111110001001, 25'b0000000000000110001110010, 25'b1111111111111001101000011, 25'b1111111111111011010001110, 25'b0000000000000101100111001, 25'b0000000000000000100100110}, 
{25'b0000000000000110111001010, 25'b0000000000000011001110001, 25'b0000000000000000000000110, 25'b1111111111111101011101001, 25'b1111111111111110101111101, 25'b1111111111111111111111001, 25'b0000000000000000000000000, 25'b1111111111111110111001001, 25'b1111111111111110000000110, 25'b1111111111111110000110101, 25'b0000000000000000000000010, 25'b0000000000000010100010001, 25'b0000000000000000000110100, 25'b0000000000000000110110001, 25'b1111111111111111010010010, 25'b0000000000000000000101111, 25'b1111111111111101100010111, 25'b0000000000000000000000100, 25'b1111111111111111101101111, 25'b1111111111111111111111011, 25'b0000000000000000000010011, 25'b0000000000000000111100110, 25'b0000000000000001100011100, 25'b0000000000000000000000000, 25'b0000000000000000000000010, 25'b1111111111110110001110110, 25'b1111111111111100110011111, 25'b0000000000000000000110110, 25'b0000000000000000010100111, 25'b0000000000000000000001010, 25'b1111111111111101001010101, 25'b0000000000000000010101111}, 
{25'b0000000000000011000000001, 25'b1111111111101111010010011, 25'b1111111111111111111111111, 25'b1111111111111110110010111, 25'b1111111111111100010001100, 25'b1111111111111111110110001, 25'b0000000000000000000000000, 25'b0000000000001000110000111, 25'b1111111111111111010011001, 25'b1111111111111111101001100, 25'b0000000000000001010100011, 25'b1111111111110101011011011, 25'b0000000000000000011000100, 25'b1111111111111000111111000, 25'b0000000000001011100011110, 25'b1111111111111111001010011, 25'b1111111111111100011000000, 25'b1111111111110111001111110, 25'b1111111111111111110101001, 25'b1111111111110100101011001, 25'b1111111111110011000010111, 25'b1111111111111111111111101, 25'b0000000000000000000000011, 25'b0000000000000000000000000, 25'b0000000000000011111001111, 25'b1111111111111111110001101, 25'b1111111111111011001110101, 25'b1111111111111110110101100, 25'b1111111111111111101000001, 25'b0000000000000000000000001, 25'b1111111111111111011111100, 25'b1111111111110100110011010}
};

localparam logic signed [24:0] bias [32] = '{
25'b0000000000000100001110011,  // 0.5280959606170654
25'b0000000000000110101110110,  // 0.8414360880851746
25'b0000000000000011001011101,  // 0.397830605506897
25'b0000000000000011010010001,  // 0.4105983078479767
25'b1111111111100010101111001,  // -3.657735586166382
25'b1111111111111000110100010,  // -0.8977976441383362
25'b0000000000001101101001000,  // 1.7051936388015747
25'b1111111111110101110010011,  // -1.2765135765075684
25'b1111111111111011010101000,  // -0.5837795734405518
25'b0000000000010101100110001,  // 2.699671983718872
25'b0000000000000001101111001,  // 0.2170683741569519
25'b0000000000000111000011010,  // 0.8814588785171509
25'b1111111111101010111011001,  // -2.634300947189331
25'b1111111111110000111110110,  // -1.877297282218933
25'b0000000000001101010011001,  // 1.6625694036483765
25'b0000000000010101111101111,  // 2.7459704875946045
25'b1111111111111100001011000,  // -0.47838035225868225
25'b0000000000001101100101101,  // 1.6984987258911133
25'b0000000000000110110101101,  // 0.8548859357833862
25'b0000000000001000000010010,  // 1.0045719146728516
25'b0000000000001011010110111,  // 1.4197649955749512
25'b0000000000000110101010001,  // 0.832463800907135
25'b0000000000000100010110001,  // 0.5434179306030273
25'b0000000000000111011010111,  // 0.9277304410934448
25'b1111111111111101010000100,  // -0.3426123857498169
25'b1111111111111011100001111,  // -0.5587119460105896
25'b1111111111111011000010000,  // -0.6208624839782715
25'b1111111111110101110000100,  // -1.2802538871765137
25'b0000000000000000011110011,  // 0.05940237268805504
25'b1111111111111001011011011,  // -0.8213341236114502
25'b0000000000000111000001101,  // 0.8783953189849854
25'b1111111111111000011001110   // -0.949700653553009
};
endpackage