// Width: 24
// NFRAC: 12
package dense_2_24_12;

localparam logic signed [23:0] weights [64][32] = '{ 
{24'b000000000000010001001101, 24'b000000000000000000100001, 24'b111111111111110011110110, 24'b111111111111111110101001, 24'b000000000000010000101101, 24'b000000000000000000000000, 24'b111111111111110110110000, 24'b111111111111111111111111, 24'b111111111111101110011110, 24'b000000000000000101000110, 24'b000000000000000000000000, 24'b111111111111111111101000, 24'b111111111111111111111110, 24'b111111111111110011001100, 24'b111111111111111100110000, 24'b111111111111101111001111, 24'b000000000000000000000000, 24'b111111111111111111001010, 24'b111111111111110011110011, 24'b111111111111110101110111, 24'b000000000000000000000000, 24'b000000000000000000000000, 24'b111111111111111111011111, 24'b111111111111111111110100, 24'b000000000000000000000000, 24'b000000000000000110011011, 24'b000000000000011000101101, 24'b000000000000001011001101, 24'b111111111111111111111110, 24'b000000000000000011001111, 24'b111111111111100101110011, 24'b000000000000000000000001}, 
{24'b111111111111111001100101, 24'b111111111111110110000101, 24'b111111111111110111001001, 24'b111111111111111100011100, 24'b111111111111111111101000, 24'b000000000000000010110000, 24'b111111111111110001101101, 24'b000000000000000000010101, 24'b000000000000000000010011, 24'b111111111111111011111110, 24'b000000000000001001111111, 24'b111111111111111101001110, 24'b111111111111111100001110, 24'b111111111111110010000111, 24'b000000000000000000011110, 24'b111111111111111100111011, 24'b000000000000000000110011, 24'b111111111111110011100010, 24'b000000000000001010111111, 24'b000000000000001110101100, 24'b111111111111111101111111, 24'b111111111111111111101000, 24'b111111111111111111111110, 24'b000000000000000001100000, 24'b111111111111111011011100, 24'b000000000000010001100110, 24'b000000000000001111110110, 24'b000000000000000000100010, 24'b000000000000000001110100, 24'b111111111111100000110110, 24'b000000000000000000011110, 24'b000000000000000000000000}, 
{24'b000000000000000100101000, 24'b111111111111111000101010, 24'b111111111111110111101101, 24'b111111111111111101010100, 24'b111111111111111011000010, 24'b111111111111111010100010, 24'b111111111111110100001010, 24'b000000000000000000010010, 24'b111111111111110111010111, 24'b000000000000000000100100, 24'b000000000000000000001000, 24'b111111111111111010110101, 24'b000000000000000101110010, 24'b111111111111111011110111, 24'b111111111111111111111010, 24'b111111111111111101101001, 24'b000000000000000000010100, 24'b000000000000000110000111, 24'b000000000000000011110000, 24'b000000000000001110101101, 24'b000000000000000010101000, 24'b111111111111111010100111, 24'b000000000000000000000001, 24'b000000000000000010001111, 24'b111111111111111110110100, 24'b000000000000001101011001, 24'b000000000000001001100011, 24'b000000000000000110001100, 24'b111111111111111111111110, 24'b111111111111110110010001, 24'b111111111111111111001000, 24'b000000000000000110010110}, 
{24'b000000000000001000110101, 24'b000000000000000001001110, 24'b000000000000000011011000, 24'b111111111111111111011000, 24'b111111111111011111011010, 24'b000000000000000000000000, 24'b000000000000000000000001, 24'b000000000000001110011110, 24'b000000000000001111100001, 24'b111111111111111111001001, 24'b111111111111111111111111, 24'b000000000000000000000000, 24'b000000000000000000000001, 24'b000000000000000000010100, 24'b111111111111111110110101, 24'b000000000000001101101111, 24'b000000000000000000000000, 24'b111111111111111110011011, 24'b111111111111111111111111, 24'b111111111111110100101110, 24'b111111111111111100000101, 24'b000000000000000011001010, 24'b111111111111111011111100, 24'b111111111111111111111110, 24'b000000000000000000001111, 24'b111111111111111100110000, 24'b000000000000000100101011, 24'b111111111111111111111111, 24'b111111111111111111111111, 24'b111111111111111111111111, 24'b111111111111110010001110, 24'b000000000000010011110110}, 
{24'b111111111111010100010100, 24'b111111111111111110011010, 24'b111111111111111111101110, 24'b000000000000000000010101, 24'b111111111111111110010100, 24'b000000000000000000011011, 24'b111111111111111100110110, 24'b111111111111110110011010, 24'b000000000000000011011110, 24'b111111111111111110101101, 24'b111111111111111111001000, 24'b111111111111111111111111, 24'b111111111111111111111111, 24'b000000000000001101011101, 24'b000000000000000000000000, 24'b000000000000010101000011, 24'b111111111111111111111111, 24'b000000000000001101111101, 24'b111111111111100110011001, 24'b000000000000000000000001, 24'b111111111111111000110110, 24'b000000000000001010110010, 24'b000000000000010000100001, 24'b000000000000000000000000, 24'b000000000000000010111001, 24'b000000000000001010011011, 24'b000000000000001111010001, 24'b000000000000000001000111, 24'b111111111111111111101101, 24'b111111111111111111111111, 24'b111111111111111111000111, 24'b000000000000001110011110}, 
{24'b000000000000000011101100, 24'b111111111111111111111111, 24'b000000000000001001100011, 24'b111111111111010110011111, 24'b111111111110100111110111, 24'b111111111111101001100100, 24'b000000000000010110101010, 24'b111111111111011000001011, 24'b111111111111111111111110, 24'b111111111111010100101001, 24'b111111111111011111111011, 24'b111111111111101010001011, 24'b000000000000010110100111, 24'b111111111111111111111111, 24'b111111111111111111000011, 24'b000000000000000000000000, 24'b111111111111111111111111, 24'b111111111111111111111110, 24'b111111111111110111100010, 24'b111111111111111111111111, 24'b111111111111100000101100, 24'b000000000000000000000000, 24'b000000000000001011111001, 24'b111111111111111111111111, 24'b000000000000000001011010, 24'b000000000000010001001000, 24'b000000000000000011010001, 24'b111111111111111111111111, 24'b111111111111111111111111, 24'b000000000000001101001010, 24'b111111111111111101110100, 24'b000000000000001100110101}, 
{24'b111111111111111101101100, 24'b111111111111110101111011, 24'b111111111111110000100010, 24'b111111111111111100111111, 24'b111111111111101101100010, 24'b000000000000000100001110, 24'b111111111111110100011110, 24'b111111111111110110111010, 24'b111111111111100101011101, 24'b000000000000000011000110, 24'b111111111111111111101011, 24'b111111111111110101110100, 24'b000000000000000111100111, 24'b111111111111111111010110, 24'b111111111111111101010110, 24'b111111111111011100100100, 24'b111111111111111111111111, 24'b000000000000000101011000, 24'b000000000000001100010001, 24'b111111111111110101100111, 24'b111111111111110110011001, 24'b111111111111111011111111, 24'b111111111111111111111010, 24'b000000000000000001110001, 24'b111111111111111101000101, 24'b111111111111010110100001, 24'b111111111111101111000010, 24'b111111111111111101000111, 24'b000000000000000000010111, 24'b111111111111111110101000, 24'b000000000000000001111101, 24'b111111111111111111111101}, 
{24'b111111111111110110001011, 24'b111111111111111010001101, 24'b111111111111111010111010, 24'b111111111111110000110100, 24'b111111111111111000100101, 24'b111111111111111111111110, 24'b000000000000000110101011, 24'b111111111111111010111100, 24'b000000000000001100110101, 24'b000000000000000000000000, 24'b000000000000000000000000, 24'b111111111111111111111111, 24'b000000000000001110000000, 24'b000000000000000000000000, 24'b111111111111111111111111, 24'b111111111111111011011110, 24'b111111111111111111111110, 24'b000000000000000000000000, 24'b111111111111111111111110, 24'b000000000000000000000000, 24'b111111111111111111111110, 24'b111111111111111111111101, 24'b000000000000000000000000, 24'b111111111111111111111111, 24'b000000000000000010110100, 24'b111111111111110100011110, 24'b000000000000000000111000, 24'b111111111111111111111110, 24'b111111111111111011011000, 24'b111111111111111111111101, 24'b000000000000000000000001, 24'b111111111111111111111111}, 
{24'b111111111111100001011100, 24'b111111111111111100010110, 24'b111111111111100111101011, 24'b000000000000000111110100, 24'b000000000000011111001010, 24'b111111111111111111111111, 24'b111111111111111110001001, 24'b000000000000001111010010, 24'b111111111111100011111010, 24'b111111111111111101000000, 24'b000000000000000000000000, 24'b111111111111110011000110, 24'b111111111111111111111110, 24'b000000000000000100110111, 24'b111111111111110011110011, 24'b000000000000110000010000, 24'b111111111111111111011100, 24'b000000000000000010111111, 24'b000000000000001101010010, 24'b000000000000001111101011, 24'b000000000000000000000000, 24'b111111111111101010100000, 24'b000000000000000000000000, 24'b000000000000011010010101, 24'b111111111111110100011001, 24'b000000000000101100101001, 24'b111111111111110110011100, 24'b111111111111110010111100, 24'b111111111111100001110010, 24'b111111111111100010010010, 24'b000000000000000000000001, 24'b000000000000000011011010}, 
{24'b000000000000000000000000, 24'b111111111111111111000000, 24'b111111111111111011010001, 24'b000000000000000000000000, 24'b000000000000010011101111, 24'b111111111111111110101101, 24'b111111111111111011111011, 24'b000000000000000101111000, 24'b000000000000000110011111, 24'b000000000000000000001110, 24'b111111111111111111011101, 24'b111111111111111111111110, 24'b111111111111111111111111, 24'b111111111111111000101110, 24'b111111111111111111111111, 24'b000000000000000000000001, 24'b000000000000000000000000, 24'b111111111111111111101011, 24'b000000000000000000001000, 24'b000000000000000101011011, 24'b000000000000000001001110, 24'b111111111111111111111111, 24'b000000000000000000000000, 24'b000000000000000000011101, 24'b000000000000000010011101, 24'b111111111111110111100011, 24'b000000000000000100010110, 24'b000000000000001111111010, 24'b111111111111111111111111, 24'b000000000000000000011001, 24'b000000000000000011001011, 24'b000000000000000100011100}, 
{24'b000000000000000110001010, 24'b000000000000000000000000, 24'b111111111111111001011001, 24'b111111111111101111111100, 24'b111111111111001101001011, 24'b000000000000001000100001, 24'b000000000000000000000001, 24'b111111111111001011000011, 24'b000000000000000010010100, 24'b111111111111111111111110, 24'b000000000000000000001111, 24'b111111111111111111111001, 24'b000000000000000000101011, 24'b000000000000000000000000, 24'b111111111111111110110010, 24'b111111111111100111100100, 24'b111111111111111111111111, 24'b000000000000001110000100, 24'b000000000000001000000101, 24'b000000000000001100001111, 24'b111111111111100011110111, 24'b111111111111101001001110, 24'b000000000000000111101011, 24'b111111111111111101110001, 24'b111111111111111101000011, 24'b000000000000010110111100, 24'b111111111111111001110100, 24'b111111111111111111111110, 24'b111111111111111111111111, 24'b000000000000001101100000, 24'b111111111111111111111111, 24'b000000000000000000011001}, 
{24'b111111111111110011010111, 24'b111111111111100000011100, 24'b000000000000000000000000, 24'b111111111111111111110111, 24'b000000000000010101010000, 24'b111111111111101110110001, 24'b111111111111110001110101, 24'b000000000000000111011010, 24'b111111111111111111111101, 24'b000000000000001001100001, 24'b000000000000000100101111, 24'b111111111111111011001010, 24'b000000000000000000000001, 24'b000000000000000000111001, 24'b111111111111111110101001, 24'b111111111111101111110011, 24'b000000000000001011001110, 24'b000000000000000001110100, 24'b000000000000010011000001, 24'b000000000000000101100010, 24'b000000000000000000000000, 24'b111111111111111101100101, 24'b000000000000001000000100, 24'b111111111111111010011110, 24'b111111111111101100010010, 24'b111111111111111111100100, 24'b000000000000001011110101, 24'b111111111111111111111111, 24'b000000000000000000100010, 24'b111111111111111001111100, 24'b000000000000001000110011, 24'b000000000000010001101011}, 
{24'b000000000000000000111110, 24'b000000000000000000000000, 24'b000000000000001110000010, 24'b000000000000000000100010, 24'b111111111111111101011001, 24'b000000000000001011100011, 24'b000000000000000101111001, 24'b111111111111111111111110, 24'b000000000000000000000011, 24'b111111111111110111000001, 24'b111111111111111100100000, 24'b111111111111110101010010, 24'b111111111111111111111111, 24'b000000000000000011001110, 24'b111111111111111011100101, 24'b000000000000110101111101, 24'b000000000000000000000001, 24'b111111111111111001111110, 24'b111111111111110011111011, 24'b111111111111111111001001, 24'b000000000000001100101101, 24'b000000000000001000001100, 24'b000000000000000000000000, 24'b111111111111111111110101, 24'b000000000000001110000011, 24'b000000000000010001001010, 24'b000000000000011111101100, 24'b000000000000000000101010, 24'b000000000000000000000000, 24'b000000000000000000000001, 24'b111111111111111111001111, 24'b111111111111111011011011}, 
{24'b111111111111110110000000, 24'b000000000000000011000110, 24'b000000000000000010100001, 24'b111111111111110000001011, 24'b111111111111101110110000, 24'b000000000000011110000000, 24'b000000000000000011001001, 24'b000000000000000000000000, 24'b111111111111110101101101, 24'b111111111111111010010110, 24'b000000000000001000010010, 24'b000000000000000100100010, 24'b000000000000000000000010, 24'b111111111111111010111110, 24'b000000000000010010010011, 24'b111111111111111111111111, 24'b111111111111111111001000, 24'b000000000000000000000000, 24'b000000000000000000110101, 24'b111111111111111101000001, 24'b000000000000000101000000, 24'b000000000000000001000000, 24'b000000000000000111010011, 24'b111111111111111111111110, 24'b000000000000000000001101, 24'b000000000000101010000111, 24'b111111111111111100011001, 24'b111111111111111110100001, 24'b111111111111111111111111, 24'b111111111111111001000000, 24'b111111111111111101011011, 24'b000000000000001011010000}, 
{24'b000000000000000011110001, 24'b000000000000000100101111, 24'b000000000000010100111001, 24'b111111111111111101011101, 24'b000000000000000110011101, 24'b000000000000010110011101, 24'b000000000000000000000010, 24'b111111111111111110000111, 24'b000000000000000111100011, 24'b111111111111111000101101, 24'b111111111111111111111111, 24'b111111111111111000010111, 24'b000000000000000000000001, 24'b000000000000011001001010, 24'b111111111111111110110111, 24'b000000000000000000000110, 24'b000000000000001111000111, 24'b000000000000000000000010, 24'b000000000000000000001100, 24'b111111111111101011111110, 24'b111111111111110000010010, 24'b111111111111111101101100, 24'b111111111111111111111111, 24'b111111111111110110101010, 24'b111111111111111101101100, 24'b111111111111111010101110, 24'b111111111111110011011011, 24'b111111111111110010011001, 24'b000000000000000001111011, 24'b000000000000000111001001, 24'b111111111111100110100100, 24'b000000000000000000001101}, 
{24'b111111111111101100111001, 24'b000000000000000000000000, 24'b111111111111111111000011, 24'b111111111111111100110100, 24'b111111111111111111111111, 24'b000000000000001000100010, 24'b111111111111111011000011, 24'b000000000000010001010110, 24'b111111111111101000110000, 24'b111111111111111111111101, 24'b000000000000000000000000, 24'b111111111111111111111111, 24'b000000000000000000000001, 24'b000000000000000000000000, 24'b111111111111111111110000, 24'b111111111111111010001100, 24'b000000000000000101000100, 24'b000000000000001011101110, 24'b111111111111111111011001, 24'b111111111111101111111010, 24'b111111111111111100001111, 24'b000000000000000111001010, 24'b000000000000000100000010, 24'b000000000000000000000001, 24'b000000000000000000001100, 24'b000000000000000101001110, 24'b111111111111110000101011, 24'b000000000000000000000000, 24'b111111111111111111111111, 24'b000000000000000000001101, 24'b000000000000000000000010, 24'b111111111111110111111100}, 
{24'b111111111111101010011111, 24'b111111111111111111101000, 24'b111111111111111111110011, 24'b111111111111111110111000, 24'b111111111111111111101100, 24'b000000000000000110110000, 24'b000000000000000000011011, 24'b000000000000000010001101, 24'b000000000000000010011100, 24'b000000000000000100000001, 24'b000000000000000101000011, 24'b000000000000001010010100, 24'b000000000000000001101101, 24'b111111111111111001110011, 24'b000000000000000000000010, 24'b000000000000011000011010, 24'b000000000000000000000001, 24'b000000000000000000000100, 24'b111111111111111111110101, 24'b000000000000000111000010, 24'b000000000000001001000111, 24'b000000000000000001111110, 24'b000000000000000010101000, 24'b111111111111111110000110, 24'b111111111111111101111100, 24'b000000000000000001101100, 24'b111111111111111011101101, 24'b111111111111110111111001, 24'b000000000000001101011010, 24'b111111111111111110000010, 24'b000000000000000010000001, 24'b111111111111110011111110}, 
{24'b000000000000000000000000, 24'b111111111111111111111111, 24'b000000000000000010011010, 24'b000000000000000000000000, 24'b000000000000111010000001, 24'b111111111111111111111100, 24'b000000000000000000000000, 24'b111111111111111111111111, 24'b000000000000000111000001, 24'b111111111111111011001100, 24'b000000000000000000000000, 24'b000000000000000000000000, 24'b000000000000000000000100, 24'b000000000000001000010000, 24'b000000000000000000000000, 24'b111111111111110110101100, 24'b111111111111111111111111, 24'b111111111111111011101101, 24'b000000000000010100111101, 24'b000000000000000000000000, 24'b111111111111111111111111, 24'b111111111111111111111110, 24'b000000000000000000000000, 24'b111111111111111111111111, 24'b000000000000000000000000, 24'b000000000000000100010111, 24'b000000000000000000000000, 24'b000000000000000000000000, 24'b111111111111111111111111, 24'b111111111111111111111111, 24'b000000000000000000000000, 24'b000000000000000010101001}, 
{24'b111111111111111111110010, 24'b000000000000000001110110, 24'b111111111111111111111100, 24'b000000000000000011000100, 24'b111111111111111101001010, 24'b111111111111111000010111, 24'b111111111111111100000000, 24'b000000000000010001110001, 24'b000000000000000000000001, 24'b000000000000000110001100, 24'b111111111111111111010010, 24'b000000000000000100001001, 24'b111111111111111101111000, 24'b111111111111110101111010, 24'b111111111111110011110011, 24'b000000000000000000110101, 24'b111111111111111111111111, 24'b111111111111111101110001, 24'b000000000000000000000000, 24'b000000000000000000000001, 24'b111111111111111111111101, 24'b000000000000000100110110, 24'b000000000000000010010010, 24'b111111111111110111111100, 24'b000000000000000111001001, 24'b111111111111110101011110, 24'b000000000000000000001000, 24'b000000000000000000000000, 24'b111111111111110101010001, 24'b000000000000000000000000, 24'b000000000000000010111010, 24'b111111111111111110000000}, 
{24'b111111111111111111010000, 24'b111111111111111001101010, 24'b000000000000000000000000, 24'b111111111111111100001011, 24'b000000000000001101110100, 24'b111111111111111111111110, 24'b111111111111111110101010, 24'b000000000000000110110101, 24'b111111111111100110111111, 24'b000000000000000000000000, 24'b111111111111111101100010, 24'b111111111111111111110111, 24'b000000000000010110011111, 24'b000000000000001110101011, 24'b111111111111111001101001, 24'b111111111111111110101010, 24'b111111111111111111111110, 24'b000000000000000000000010, 24'b111111111111111111111111, 24'b000000000000000000000001, 24'b000000000000000000000000, 24'b111111111111110111010011, 24'b111111111111111000011000, 24'b000000000000001000011000, 24'b000000000000000000000000, 24'b111111111111110111001110, 24'b000000000000000001100100, 24'b111111111111111010110110, 24'b111111111111111101110111, 24'b000000000000001000101100, 24'b000000000000000000000010, 24'b111111111111110000001011}, 
{24'b000000000000101000100111, 24'b000000000000010101111000, 24'b111111111111110000000010, 24'b000000000000000000001101, 24'b111111111111101001110110, 24'b000000000000000000000000, 24'b000000000000001110010000, 24'b000000000000000001111111, 24'b000000000000001110010100, 24'b111111111111111111111110, 24'b111111111111110110000101, 24'b111111111111111010111110, 24'b000000000000001001000100, 24'b000000000000000001110001, 24'b111111111111111001101101, 24'b000000000000001000011011, 24'b000000000000100010010000, 24'b111111111111110111101011, 24'b111111111111101101000011, 24'b000000000000000000000000, 24'b111111111111111110001010, 24'b111111111111110100101100, 24'b111111111111111111001110, 24'b111111111111111111111001, 24'b000000000000000101100000, 24'b111111111111101000111011, 24'b000000000000000101101100, 24'b111111111111111111111011, 24'b000000000000000000000001, 24'b000000000000000110111110, 24'b111111111111111110001001, 24'b000000000000000011110100}, 
{24'b111111111111111010000100, 24'b111111111111110011101101, 24'b111111111111111101101011, 24'b111111111111110101010010, 24'b111111111111111110111001, 24'b000000000000000011001001, 24'b000000000000000000000000, 24'b111111111111111111010001, 24'b000000000000000010011010, 24'b111111111111111111110001, 24'b000000000000000000000000, 24'b111111111111110010000111, 24'b000000000000000110100001, 24'b000000000000000101001001, 24'b111111111111111001011100, 24'b000000000000011100011000, 24'b111111111111111111111111, 24'b000000000000000000000000, 24'b111111111111111111101111, 24'b000000000000000000000000, 24'b000000000000010100001110, 24'b111111111111100001111000, 24'b111111111111111001000100, 24'b111111111111111100011010, 24'b111111111111111110110011, 24'b000000000000001100100111, 24'b111111111111111100101001, 24'b000000000000000001001000, 24'b000000000000011110111111, 24'b111111111111011111001100, 24'b111111111111101000100000, 24'b000000000000000001011011}, 
{24'b000000000000000001000100, 24'b111111111111111100001111, 24'b111111111111111111111111, 24'b000000000000000000000000, 24'b111111111111010001111111, 24'b111111111111011001001100, 24'b000000000000000000000110, 24'b111111111111111111111111, 24'b111111111111101111000010, 24'b000000000000000001100101, 24'b000000000000000000000000, 24'b111111111111111110001111, 24'b000000000000000000000000, 24'b111111111111111100010000, 24'b111111111111111100101000, 24'b111111111111111011100101, 24'b111111111111110110100101, 24'b000000000000010010000100, 24'b000000000000000000000000, 24'b000000000000000010111101, 24'b111111111111111111111110, 24'b111111111111111011011111, 24'b000000000000000000000000, 24'b111111111111111010011100, 24'b000000000000001110000011, 24'b111111111111011000001010, 24'b000000000000001110000101, 24'b111111111111111111111111, 24'b111111111111111111101100, 24'b000000000000001100110011, 24'b111111111111111111111111, 24'b000000000000001111000111}, 
{24'b111111111111111111111111, 24'b000000000000000000010101, 24'b111111111111111101001111, 24'b000000000000000100110011, 24'b000000000000000011100010, 24'b111111111111101010000111, 24'b000000000000000000000000, 24'b000000000000000100000111, 24'b000000000000100101000110, 24'b111111111111111111011011, 24'b000000000000000000000000, 24'b000000000000000011100110, 24'b000000000000010110111110, 24'b111111111111111101111101, 24'b000000000000000000111001, 24'b000000000000000110011101, 24'b111111111111111111111111, 24'b000000000000000001110001, 24'b111111111111111111111110, 24'b000000000000000000000011, 24'b111111111111101110011110, 24'b000000000000000010011101, 24'b000000000000000100011111, 24'b000000000000000001011101, 24'b111111111111111111111111, 24'b000000000000001101111110, 24'b000000000000000000010010, 24'b000000000000001000000100, 24'b111111111111100101010001, 24'b000000000000000110100101, 24'b000000000000011001010100, 24'b000000000000000000010111}, 
{24'b111111111111101001100010, 24'b000000000000001101100000, 24'b111111111111101111010101, 24'b000000000000000111110111, 24'b111111111111111001010000, 24'b000000000000000000000001, 24'b000000000000011111110110, 24'b111111111111110001000110, 24'b111111111111101101010111, 24'b000000000000001010111101, 24'b111111111111110001101111, 24'b111111111111111110011111, 24'b111111111111111111111100, 24'b000000000000010110000001, 24'b111111111111111111111001, 24'b111111111111101100101100, 24'b111111111111111111111111, 24'b000000000000011100001101, 24'b111111111111100001110110, 24'b111111111111111110011100, 24'b000000000000010100010000, 24'b111111111111101000110010, 24'b000000000000000011011001, 24'b111111111111111111000010, 24'b000000000000010001010111, 24'b111111111111011111011100, 24'b111111111111101000110010, 24'b111111111111110011011100, 24'b111111111111111111111111, 24'b000000000000000110101000, 24'b000000000000000001100110, 24'b000000000000001011011010}, 
{24'b111111111111111010001100, 24'b000000000000000011010100, 24'b111111111111111111111111, 24'b000000000000001001100101, 24'b111111111111111101100100, 24'b000000000000001110100001, 24'b000000000000000000001000, 24'b111111111111111111010010, 24'b111111111111111111110111, 24'b000000000000000000000100, 24'b000000000000000000000000, 24'b111111111111111111111111, 24'b111111111111111111111000, 24'b000000000000100001010010, 24'b000000000000000000110011, 24'b000000000000001100000101, 24'b000000000000000000000001, 24'b111111111111110010011101, 24'b111111111111111011000111, 24'b111111111111111111111111, 24'b111111111111111110111100, 24'b000000000000000010101100, 24'b111111111111111111111111, 24'b111111111111110100001001, 24'b111111111111111111111111, 24'b000000000000010010111010, 24'b000000000000010011110110, 24'b111111111111111111111111, 24'b111111111111111110111101, 24'b000000000000000000000000, 24'b111111111111111111111101, 24'b111111111111111001110101}, 
{24'b111111111111111010110101, 24'b000000000000000000000000, 24'b000000000000010001011110, 24'b000000000000000000000000, 24'b000000000000000000000000, 24'b111111111111111000101110, 24'b000000000000000000000001, 24'b111111111111001000101110, 24'b000000000000001101110010, 24'b000000000000000000111000, 24'b000000000000000001101101, 24'b111111111111101000111110, 24'b000000000000000000001101, 24'b111111111111110111001101, 24'b111111111111111101111000, 24'b000000000000000000000000, 24'b000000000000000001010000, 24'b000000000000000000000000, 24'b000000000000000111001100, 24'b000000000000000000000001, 24'b111111111111111111011011, 24'b000000000000010101000100, 24'b000000000000011000000110, 24'b111111111111110001110111, 24'b111111111111110110111010, 24'b000000000000001111111110, 24'b111111111111101100011100, 24'b000000000000000001111000, 24'b111111111111111111111101, 24'b111111111111111111111111, 24'b111111111111111111111111, 24'b000000000000001011110010}, 
{24'b111111111111111000101111, 24'b111111111111111111111101, 24'b111111111111110000101100, 24'b111111111111110011000100, 24'b111111111111111111000111, 24'b111111111111110111010111, 24'b000000000000000000000000, 24'b000000000000000101110101, 24'b111111111111110000101010, 24'b111111111111111010101010, 24'b111111111111111100110100, 24'b000000000000000000000001, 24'b000000000000000001110010, 24'b111111111111111111010111, 24'b111111111111111100000110, 24'b000000000000000110000111, 24'b000000000000001110010000, 24'b000000000000001000011001, 24'b111111111111110111101000, 24'b000000000000000011000111, 24'b111111111111111111001111, 24'b111111111111111110001011, 24'b000000000000000001011100, 24'b000000000000000001000001, 24'b111111111111111011100011, 24'b000000000000000101101100, 24'b111111111111111010001100, 24'b000000000000000011110101, 24'b111111111111111111111111, 24'b111111111111101101000110, 24'b111111111111111110010100, 24'b000000000000001110011001}, 
{24'b111111111111111110010001, 24'b111111111111111010101101, 24'b000000000000000100111011, 24'b000000000000010000001100, 24'b000000000000000101011011, 24'b000000000000000101010001, 24'b000000000000000010111111, 24'b111111111111110011000110, 24'b111111111111110010110111, 24'b000000000000000100011000, 24'b000000000000000000110001, 24'b000000000000000010110000, 24'b000000000000000001011011, 24'b000000000000000000010110, 24'b000000000000001101001000, 24'b000000000000000000011110, 24'b111111111111111100100011, 24'b000000000000000110100111, 24'b111111111111111110000110, 24'b111111111111111101101101, 24'b000000000000000111000010, 24'b111111111111111000000100, 24'b111111111111111110010010, 24'b000000000000001000001000, 24'b000000000000000001011010, 24'b111111111111111001001011, 24'b111111111111110011010101, 24'b111111111111111111001111, 24'b111111111111101110001000, 24'b000000000000000011110110, 24'b000000000000000110100000, 24'b000000000000000000000100}, 
{24'b111111111111111111001000, 24'b111111111111111110101111, 24'b111111111111111111001111, 24'b111111111111111101110010, 24'b111111111111110111100101, 24'b111111111111110111000001, 24'b000000000000000100000010, 24'b000000000000000000100001, 24'b111111111111110100010100, 24'b000000000000001010101101, 24'b111111111111111110101010, 24'b111111111111111111111101, 24'b111111111111111000111100, 24'b000000000000000000010101, 24'b000000000000000001111000, 24'b111111111111111100101000, 24'b111111111111111110111110, 24'b111111111111111101010101, 24'b111111111111111010110110, 24'b000000000000000000000001, 24'b111111111111110111000000, 24'b000000000000000110100001, 24'b111111111111110010011101, 24'b000000000000000000010100, 24'b000000000000000010101011, 24'b000000000000000111111011, 24'b000000000000000001101100, 24'b000000000000000000011000, 24'b000000000000010010101100, 24'b000000000000000011010011, 24'b000000000000000000000001, 24'b000000000000000101010111}, 
{24'b111111111111111110110000, 24'b000000000000010000001011, 24'b111111111111111111111111, 24'b111111111111111101111001, 24'b111111111111110010010100, 24'b111111111111111011001100, 24'b000000000000011010010101, 24'b111111111111010011111001, 24'b111111111111101001101000, 24'b111111111111110011001110, 24'b111111111111110001111101, 24'b111111111111101111110001, 24'b111111111111111111111101, 24'b000000000000011110111111, 24'b111111111111111110010100, 24'b000000000000000000000000, 24'b111111111111110010011111, 24'b000000000000011100100001, 24'b111111111111100101100101, 24'b000000000000000000000000, 24'b111111111111111111111110, 24'b111111111111101010011110, 24'b000000000000000000000000, 24'b111111111111111111111111, 24'b000000000000000011100110, 24'b111111111111111100010100, 24'b111111111111110110100010, 24'b111111111111111111111111, 24'b000000000000001011001011, 24'b000000000000000000001101, 24'b111111111111111010110111, 24'b000000000000000000000011}, 
{24'b000000000000010111100011, 24'b111111111111111000110101, 24'b000000000000001000011100, 24'b111111111111111101111011, 24'b000000000000000100111000, 24'b111111111111111111110000, 24'b111111111111111111110100, 24'b111111111111111010000011, 24'b000000000000000000000001, 24'b000000000000000101111001, 24'b111111111111111111111111, 24'b111111111111111100001111, 24'b111111111111111111111110, 24'b000000000000001110101000, 24'b000000000000000001001110, 24'b000000000000000010100101, 24'b000000000000000001100010, 24'b111111111111111110011101, 24'b000000000000000001010011, 24'b000000000000000000000000, 24'b111111111111111111011011, 24'b111111111111111111111111, 24'b111111111111101100011100, 24'b111111111111111111111111, 24'b000000000000000011101100, 24'b111111111111111000100011, 24'b111111111111110111010110, 24'b111111111111111111111111, 24'b111111111111111111111100, 24'b000000000000100011101100, 24'b111111111111101101101101, 24'b111111111111111000100100}, 
{24'b111111111111111101001011, 24'b111111111111111001011001, 24'b111111111111111011110111, 24'b000000000000000010010100, 24'b000000000000001000111011, 24'b111111111111110111101100, 24'b111111111111111111111010, 24'b111111111111110001111011, 24'b000000000000000011111000, 24'b000000000000001000101101, 24'b111111111111110010010101, 24'b111111111111101111110100, 24'b000000000000000001100001, 24'b111111111111010100010000, 24'b111111111111111011001011, 24'b111111111111111000000110, 24'b111111111111110011010101, 24'b111111111111111111111110, 24'b000000000000001000100101, 24'b000000000000000000000000, 24'b111111111111111101000101, 24'b111111111111111101001001, 24'b000000000000000000000000, 24'b000000000000000000000000, 24'b111111111111111100001110, 24'b111111111111001111101110, 24'b111111111111011100011101, 24'b111111111111101110100011, 24'b000000000000000011100101, 24'b000000000000001101001100, 24'b111111111111111111111110, 24'b000000000000001111011000}, 
{24'b111111111111111010000110, 24'b111111111111110010010000, 24'b000000000000001010011110, 24'b000000000000000100110001, 24'b000000000000000010110001, 24'b111111111111111010000111, 24'b111111111111111101111010, 24'b000000000000000110010011, 24'b000000000000100010011111, 24'b111111111111110101000010, 24'b111111111111111111111111, 24'b111111111111111111111111, 24'b000000000000000111100001, 24'b111111111111111100011111, 24'b111111111111111110110110, 24'b111111111111111110111011, 24'b111111111111111001100110, 24'b111111111111111111111100, 24'b000000000000000000000000, 24'b000000000000001110100000, 24'b111111111111110111011111, 24'b111111111111111111110011, 24'b000000000000001000001110, 24'b111111111111111111010110, 24'b000000000000000000000000, 24'b000000000000100001101011, 24'b000000000000010100110000, 24'b000000000000000000001101, 24'b000000000000000000000001, 24'b111111111111100101000100, 24'b111111111111111011101000, 24'b111111111111111111111111}, 
{24'b000000000000000000111101, 24'b000000000000000011000101, 24'b111111111111111111000111, 24'b000000000000000000000000, 24'b000000000000001110110011, 24'b111111111111100001000100, 24'b000000000000000000000000, 24'b111111111111111001111010, 24'b000000000000001011111011, 24'b000000000000000000000000, 24'b111111111111111110110100, 24'b000000000000000000000000, 24'b000000000000000000000001, 24'b111111111111111111111111, 24'b000000000000000000010111, 24'b111111111111111001000111, 24'b000000000000010000100110, 24'b111111111111111111101001, 24'b111111111111111111000000, 24'b111111111111111111111111, 24'b000000000000000000000001, 24'b111111111111111111100000, 24'b000000000000000000000001, 24'b111111111111111111111111, 24'b000000000000000000110100, 24'b111111111111101011101101, 24'b000000000000000011010011, 24'b000000000000001011101110, 24'b111111111111111111110010, 24'b000000000000000110000010, 24'b111111111111111111111110, 24'b000000000000000100110010}, 
{24'b111111111111110011000111, 24'b000000000000000000100101, 24'b111111111111100001001000, 24'b000000000000000000011100, 24'b111111111111111100110011, 24'b111111111111111101011101, 24'b111111111111111111111010, 24'b111111111111111010001010, 24'b111111111111111101101100, 24'b111111111111111011110100, 24'b000000000000000011000000, 24'b000000000000000001101110, 24'b111111111111110100101001, 24'b000000000000000000000010, 24'b111111111111111111111000, 24'b111111111111111111011110, 24'b000000000000000100100000, 24'b111111111111111110101101, 24'b111111111111111110001111, 24'b111111111111111110001001, 24'b111111111111111111111100, 24'b000000000000010001010110, 24'b111111111111111111111111, 24'b000000000000000000000000, 24'b111111111111111111011001, 24'b000000000000010100010011, 24'b000000000000001100000100, 24'b000000000000000010001011, 24'b111111111111111001110101, 24'b111111111111111111010111, 24'b000000000000000100001011, 24'b000000000000000011101011}, 
{24'b000000000000000010001011, 24'b000000000000000010100000, 24'b111111111111111111111111, 24'b000000000000000000000001, 24'b111111111111100010000000, 24'b000000000000000010110010, 24'b000000000000000001100101, 24'b111111111111111111111110, 24'b000000000000000000000010, 24'b111111111111110101001001, 24'b111111111111111111111111, 24'b000000000000000000000000, 24'b111111111111110101101101, 24'b000000000000000000000000, 24'b000000000000000000000001, 24'b000000000000000000000001, 24'b000000000000000000000000, 24'b111111111111101001001110, 24'b000000000000000000100111, 24'b111111111111111111111101, 24'b111111111111111111111110, 24'b000000000000000000000000, 24'b000000000000001000010000, 24'b111111111111111111111111, 24'b000000000000000000000000, 24'b000000000000011101001011, 24'b000000000000010101110001, 24'b000000000000000000000000, 24'b000000000000000000000000, 24'b111111111111110001000011, 24'b000000000000000000000001, 24'b111111111111111111111111}, 
{24'b000000000000000100110110, 24'b000000000000000011011000, 24'b000000000000010000001100, 24'b111111111111110000000111, 24'b000000000000001000011110, 24'b000000000000000111100110, 24'b000000000000000000011001, 24'b000000000000001100010001, 24'b000000000000000000110000, 24'b111111111111111111001110, 24'b000000000000000010011000, 24'b000000000000000000010111, 24'b111111111111111111111101, 24'b000000000000000111101110, 24'b111111111111111111101001, 24'b111111111111111101011101, 24'b000000000000000000000010, 24'b000000000000000010000010, 24'b111111111111111100111010, 24'b000000000000000110010100, 24'b000000000000000010000101, 24'b111111111111011010110110, 24'b111111111111111000101011, 24'b000000000000000101110110, 24'b111111111111111111111111, 24'b111111111111011111101011, 24'b111111111111110111111011, 24'b111111111111111110100001, 24'b111111111111111111111101, 24'b111111111111111100010110, 24'b000000000000000000000000, 24'b111111111111111101011101}, 
{24'b000000000000000000000111, 24'b111111111111111111111111, 24'b111111111111111010001001, 24'b111111111111110101001110, 24'b000000000000000010101011, 24'b000000000000000000000000, 24'b000000000000000110000110, 24'b111111111111111111101000, 24'b000000000000001111111110, 24'b111111111111111111101111, 24'b000000000000000000000000, 24'b111111111111101010000001, 24'b111111111111111111111110, 24'b000000000000001000000011, 24'b111111111111111111111111, 24'b111111111111101111010100, 24'b000000000000000000000000, 24'b111111111111111111010001, 24'b000000000000010000110100, 24'b111111111111111111111111, 24'b111111111111100100000011, 24'b111111111111111111111111, 24'b000000000000010000100000, 24'b111111111111111111111111, 24'b111111111111111111111111, 24'b000000000000001000111000, 24'b111111111111111001111111, 24'b000000000000000100011011, 24'b000000000000000000000000, 24'b111111111111110011000110, 24'b000000000000000000000000, 24'b000000000000000000001010}, 
{24'b111111111111110010001010, 24'b000000000000000000000100, 24'b000000000000000000000010, 24'b111111111111111111100111, 24'b000000000000011111101110, 24'b111111111111111000000011, 24'b111111111111111111101001, 24'b111111111111111111100010, 24'b111111111111111101001000, 24'b111111111111111100110001, 24'b000000000000000100001011, 24'b000000000000001000100000, 24'b111111111111111101101001, 24'b000000000000001111111110, 24'b000000000000000000000000, 24'b111111111111111111111110, 24'b111111111111101101110100, 24'b111111111111111111111101, 24'b000000000000000000000001, 24'b111111111111111010111001, 24'b000000000000000000001000, 24'b000000000000000010011000, 24'b000000000000000000110110, 24'b111111111111111111011010, 24'b111111111111111100101111, 24'b111111111111110011000001, 24'b111111111111101101000100, 24'b000000000000000000000001, 24'b111111111111111000110000, 24'b000000000000000010100011, 24'b111111111111111111111110, 24'b000000000000000100110101}, 
{24'b111111111111100101100011, 24'b111111111111110101111111, 24'b111111111111110110000000, 24'b000000000000000000000000, 24'b000000000000100100100011, 24'b111111111111110001110000, 24'b000000000000000000000000, 24'b111111111111111100100010, 24'b111111111111100101110001, 24'b000000000000001000110111, 24'b111111111111111111111111, 24'b000000000000100100010011, 24'b000000000000000000000001, 24'b111111111111111100111101, 24'b111111111111111111111110, 24'b000000000000000010000001, 24'b111111111111111110110011, 24'b000000000000000000000001, 24'b111111111111111101000001, 24'b000000000000011111101101, 24'b000000000000000010011110, 24'b111111111111111101010101, 24'b000000000000000111000000, 24'b111111111111111111111110, 24'b111111111111111111111111, 24'b111111111111111001110001, 24'b111111111111111101000000, 24'b111111111111100010000011, 24'b111111111111110110110000, 24'b111111111111111111111111, 24'b111111111111111111111011, 24'b111111111111111100001111}, 
{24'b000000000000001110011101, 24'b111111111111001100110101, 24'b111111111111010001101000, 24'b111111111111110101000111, 24'b000000000000101010110101, 24'b111111111111111111111111, 24'b111111111111101001110100, 24'b000000000000010000111100, 24'b000000000000000011110011, 24'b000000000000000000000011, 24'b000000000000001101010101, 24'b111111111111101110101000, 24'b000000000000000000000011, 24'b000000000000000000010001, 24'b111111111111111101111111, 24'b000000000000000001001001, 24'b111111111111111001010110, 24'b111111111111000101000001, 24'b000000000000001010101111, 24'b000000000000010110000100, 24'b000000000000010000111101, 24'b000000000000000000001010, 24'b000000000000000001110111, 24'b111111111111100110001101, 24'b111111111111010111100000, 24'b111111111111111111101011, 24'b111111111111101100110100, 24'b111111111111100010101100, 24'b111111111111110011100001, 24'b111111111111000111110111, 24'b000000000000011010110101, 24'b000000000000011011011110}, 
{24'b000000000000000000000001, 24'b000000000000000000000010, 24'b000000000000000000001001, 24'b000000000000000000000000, 24'b000000000000010000100100, 24'b111111111111110100000010, 24'b000000000000000001001000, 24'b000000000000000100101010, 24'b111111111111101001101010, 24'b000000000000000010010110, 24'b111111111111111111101101, 24'b111111111111111111111100, 24'b111111111111111111111111, 24'b000000000000001111010101, 24'b000000000000000011010100, 24'b000000000000000001011001, 24'b000000000000000011111101, 24'b000000000000010101010101, 24'b111111111111110010000001, 24'b000000000000000000000000, 24'b111111111111110101011111, 24'b111111111111111111111110, 24'b000000000000010100001000, 24'b000000000000000000100001, 24'b111111111111111111110100, 24'b111111111111011100000101, 24'b111111111111111111011010, 24'b111111111111110110000111, 24'b111111111111111100000110, 24'b000000000000000000001110, 24'b000000000000001000101001, 24'b000000000000000110101000}, 
{24'b111111111111111101001110, 24'b000000000000001000100100, 24'b111111111111101100100011, 24'b000000000000000001010100, 24'b000000000000001100011001, 24'b111111111111111101011110, 24'b111111111111111111101101, 24'b000000000000001010011100, 24'b000000000000000000000001, 24'b111111111111111111111111, 24'b111111111111111011110100, 24'b000000000000000000000000, 24'b000000000000000000000001, 24'b111111111111111101110011, 24'b111111111111111000001101, 24'b111111111111111011110000, 24'b111111111111111100011001, 24'b111111111111111011111110, 24'b111111111111111000111110, 24'b000000000000000000000000, 24'b111111111111111111111110, 24'b111111111111111101001000, 24'b111111111111111011101111, 24'b000000000000011001011101, 24'b000000000000000000000000, 24'b111111111111101000111101, 24'b111111111111111111011101, 24'b000000000000000111111000, 24'b000000000000000000000001, 24'b000000000000000000000000, 24'b000000000000010000000011, 24'b111111111111111111111110}, 
{24'b111111111111111111111111, 24'b000000000000000000010000, 24'b111111111111111111111110, 24'b111111111111110110000000, 24'b111111111111001000111100, 24'b000000000000000000000011, 24'b000000000000000000000001, 24'b111111111111111111100101, 24'b111111111111011001101000, 24'b000000000000000101001110, 24'b111111111111111001101110, 24'b111111111111111111111111, 24'b000000000000000000000001, 24'b111111111111101000010100, 24'b111111111111111101000100, 24'b111111111111111111111110, 24'b000000000000000000000101, 24'b000000000000000000100001, 24'b000000000000000010010100, 24'b000000000000010110000110, 24'b111111111111111000010110, 24'b111111111111101100110111, 24'b000000000000000000000000, 24'b111111111111101111011111, 24'b111111111111111001101011, 24'b111111111111110001001100, 24'b111111111111111111100001, 24'b111111111111111111001100, 24'b111111111111111110110101, 24'b111111111111100001110110, 24'b111111111111111101110100, 24'b000000000000001111100000}, 
{24'b000000000000000111001111, 24'b000000000000001110000001, 24'b111111111111111111110111, 24'b000000000000001010001100, 24'b111111111111110010100000, 24'b111111111111111000000010, 24'b000000000000000110000111, 24'b000000000000000100011001, 24'b111111111111111100111111, 24'b111111111111111111111111, 24'b111111111111111111111111, 24'b111111111111111111111111, 24'b111111111111111111111110, 24'b111111111111101011011111, 24'b111111111111111111111111, 24'b000000000000001001001110, 24'b111111111111111000101011, 24'b000000000000000010001110, 24'b111111111111111111111010, 24'b111111111111111111111011, 24'b000000000000001101010001, 24'b111111111111101011000100, 24'b000000000000010001111110, 24'b000000000000000011000010, 24'b000000000000000000000001, 24'b000000000000001101100011, 24'b000000000000000000001100, 24'b111111111111111101101100, 24'b111111111111100111101001, 24'b111111111111111000111111, 24'b111111111111110101000110, 24'b000000000000001011010111}, 
{24'b000000000000000000000000, 24'b000000000000000000011101, 24'b111111111111101000100101, 24'b111111111111111111110110, 24'b000000000000001101001110, 24'b111111111111110110111100, 24'b111111111111111111001110, 24'b111111111111111111111111, 24'b000000000000000001010011, 24'b000000000000000000000000, 24'b000000000000000000000000, 24'b111111111111110010111101, 24'b000000000000000110001001, 24'b000000000000000000011000, 24'b000000000000000000000000, 24'b000000000000000010011001, 24'b111111111111111111111110, 24'b111111111111110110011110, 24'b000000000000000001001001, 24'b000000000000000000000000, 24'b111111111111111101110011, 24'b111111111111111110100110, 24'b000000000000010010111101, 24'b111111111111111111111111, 24'b000000000000000000000000, 24'b111111111111101101010001, 24'b111111111111101011000101, 24'b000000000000001111011100, 24'b111111111111111111111010, 24'b111111111111111111111110, 24'b000000000000000001110001, 24'b000000000000010010000101}, 
{24'b111111111111101010001100, 24'b111111111111111111111111, 24'b111111111111110010011000, 24'b000000000000000000010001, 24'b111111111111101001011000, 24'b000000000000000000000000, 24'b111111111111111111111110, 24'b111111111111111011110100, 24'b111111111111011101111011, 24'b111111111111111110010110, 24'b000000000000000000000000, 24'b111111111111111111011110, 24'b111111111111111111111110, 24'b000000000000000000000000, 24'b111111111111111111011100, 24'b111111111111111100110100, 24'b111111111111110110100011, 24'b111111111111111001111001, 24'b000000000000000100001111, 24'b111111111111111111110110, 24'b111111111111111110011000, 24'b000000000000000000000000, 24'b000000000000010101100011, 24'b111111111111111111111111, 24'b000000000000001001100100, 24'b000000000000000101110111, 24'b111111111111110111001100, 24'b000000000000001101101001, 24'b111111111111111101000100, 24'b000000000000000000000000, 24'b111111111111111111111011, 24'b000000000000100101010000}, 
{24'b111111111111101011111001, 24'b000000000000000001111001, 24'b000000000000000011001111, 24'b111111111111111110001101, 24'b000000000000001111101000, 24'b111111111111101100101010, 24'b111111111111111111100011, 24'b000000000000010000111111, 24'b000000000000001010001100, 24'b000000000000000000100101, 24'b111111111111111111111111, 24'b111111111111111011100111, 24'b111111111111111010010001, 24'b111111111111111011110111, 24'b111111111111111100110100, 24'b000000000000000101110001, 24'b111111111111111111111111, 24'b000000000000000000100001, 24'b000000000000001001000010, 24'b000000000000000000000000, 24'b000000000000000000000000, 24'b000000000000000000111101, 24'b000000000000010000001000, 24'b000000000000000010111011, 24'b000000000000000000011011, 24'b111111111111111001000111, 24'b111111111111111111111111, 24'b000000000000000000000000, 24'b111111111111111111000110, 24'b111111111111111111001110, 24'b111111111111111111111110, 24'b000000000000000100010100}, 
{24'b111111111111111111111111, 24'b000000000000000000001111, 24'b111111111111110010011011, 24'b111111111111111011001110, 24'b000000000000010010000011, 24'b111111111111111111111110, 24'b111111111111111011000010, 24'b000000000000001111101001, 24'b111111111111111100100111, 24'b000000000000010010101010, 24'b000000000000000101011110, 24'b111111111111111000010011, 24'b000000000000000000000010, 24'b000000000000000000001110, 24'b111111111111111111000011, 24'b000000000000000001010111, 24'b111111111111111011000100, 24'b111111111111101111001001, 24'b000000000000010001110010, 24'b000000000000001001111100, 24'b000000000000101000100111, 24'b000000000000001100110110, 24'b000000000000001111111000, 24'b111111111111111111111111, 24'b000000000000000000000000, 24'b000000000000000000000000, 24'b000000000000000011101010, 24'b000000000000000101000100, 24'b111111111111100101000111, 24'b111111111111111111111111, 24'b111111111111111111101011, 24'b111111111111111111100101}, 
{24'b000000000000000000000010, 24'b111111111111111010011001, 24'b111111111111111001010111, 24'b000000000000000000000000, 24'b111111111111110000011010, 24'b000000000000000000000000, 24'b000000000000001100010000, 24'b000000000000000110111111, 24'b000000000000000011011001, 24'b111111111111111001101011, 24'b000000000000000000000000, 24'b111111111111111111111111, 24'b111111111111111111111111, 24'b111111111111111111111111, 24'b111111111111111101010001, 24'b000000000000001100111011, 24'b111111111111111111111111, 24'b111111111111111111111101, 24'b111111111111101100101001, 24'b000000000000000000000000, 24'b111111111111110011101011, 24'b111111111111111111111011, 24'b000000000000000000000000, 24'b111111111111111111101111, 24'b000000000000000000111101, 24'b000000000000000001000111, 24'b000000000000000001110010, 24'b000000000000001000110110, 24'b111111111111111011110101, 24'b111111111111111111100000, 24'b111111111111100011010010, 24'b000000000000000101000010}, 
{24'b000000000000011100010001, 24'b111111111111111111011100, 24'b000000000000000100001111, 24'b111111111111111001010011, 24'b111111111111111010100010, 24'b000000000000000010001000, 24'b000000000000001010010000, 24'b000000000000000000000000, 24'b000000000000100001101110, 24'b000000000000000000000001, 24'b111111111111111110101000, 24'b000000000000000001001101, 24'b000000000000000110000001, 24'b111111111111111111110101, 24'b000000000000000011011010, 24'b000000000000000110100111, 24'b111111111111111111101110, 24'b111111111111100011100000, 24'b111111111111111100011001, 24'b111111111111111111111001, 24'b000000000000000111011100, 24'b000000000000000000000110, 24'b111111111111111111111110, 24'b000000000000000111001100, 24'b000000000000000001001001, 24'b111111111111101111001000, 24'b111111111111111001011011, 24'b000000000000001000011101, 24'b111111111111111110001100, 24'b000000000000010000100001, 24'b111111111111111111111011, 24'b111111111111110100100011}, 
{24'b000000000000000000110101, 24'b000000000000000110100001, 24'b111111111111111111111111, 24'b111111111111111101100001, 24'b111111111111101001011010, 24'b111111111111111111111110, 24'b000000000000000010111100, 24'b111111111111111101000011, 24'b000000000000001010100011, 24'b111111111111111101110100, 24'b111111111111111111111100, 24'b111111111111111101110111, 24'b111111111111111111111111, 24'b111111111111111101101000, 24'b000000000000000000000000, 24'b000000000000010100000010, 24'b000000000000000000000000, 24'b111111111111111111111000, 24'b111111111111111111111111, 24'b111111111111111111111111, 24'b111111111111111111111111, 24'b111111111111111111111110, 24'b000000000000000010001011, 24'b000000000000001000000011, 24'b000000000000000000000000, 24'b000000000000000000010001, 24'b000000000000000010000100, 24'b111111111111111111111101, 24'b000000000000000000000000, 24'b000000000000000001010011, 24'b000000000000000000000110, 24'b000000000000000110001100}, 
{24'b111111111111101100001111, 24'b000000000000001000010101, 24'b000000000000000001001001, 24'b111111111111111001010001, 24'b111111111111100110011100, 24'b111111111111111110110101, 24'b000000000000000100010010, 24'b111111111111100110100100, 24'b000000000000100000101111, 24'b000000000000000100100101, 24'b000000000000000001000000, 24'b000000000000000110000010, 24'b000000000000000010110101, 24'b000000000000000000000010, 24'b000000000000011010000110, 24'b111111111111111010100111, 24'b000000000000000000010101, 24'b000000000000000000000000, 24'b111111111111111111100100, 24'b000000000000000000001111, 24'b111111111111100100010111, 24'b000000000000000001000101, 24'b000000000000001001110010, 24'b000000000000000010011001, 24'b000000000000000010010011, 24'b111111111111010101111111, 24'b111111111111101010001011, 24'b111111111111110000100110, 24'b000000000000000000001010, 24'b111111111111111111111000, 24'b000000000000010100110110, 24'b111111111111110010111001}, 
{24'b111111111111111111001011, 24'b111111111111110011100011, 24'b111111111111111001011000, 24'b111111111111100101110110, 24'b111111111111101111010110, 24'b000000000000010101100001, 24'b000000000000010011110101, 24'b111111111111110101000111, 24'b000000000000000010101010, 24'b111111111111111101100001, 24'b111111111111111001111111, 24'b111111111111101111111010, 24'b000000000000000110100110, 24'b111111111111101101110100, 24'b000000000000001100000101, 24'b111111111111111111111110, 24'b000000000000010101011111, 24'b111111111111111111111111, 24'b111111111111111111100000, 24'b111111111111110111010101, 24'b111111111111111101010101, 24'b111111111111111011110111, 24'b111111111111101110111111, 24'b000000000000000101010001, 24'b111111111111111111111111, 24'b111111111111111111100110, 24'b111111111111110001011001, 24'b000000000000010100001001, 24'b000000000000010001110111, 24'b111111111111111010001101, 24'b111111111111010111101001, 24'b000000000000001001001001}, 
{24'b000000000000000000000001, 24'b111111111111111110010111, 24'b111111111111111111111111, 24'b111111111111111001110001, 24'b000000000000000001110100, 24'b000000000000000000100101, 24'b000000000000000100011101, 24'b000000000000000000010111, 24'b000000000000000111100010, 24'b111111111111111111111100, 24'b000000000000000000000000, 24'b000000000000000110000110, 24'b000000000000000000000111, 24'b000000000000000000110010, 24'b111111111111110111100001, 24'b111111111111111001000110, 24'b000000000000000000000000, 24'b000000000000001011101000, 24'b000000000000000011101000, 24'b000000000000001000000011, 24'b111111111111111110111100, 24'b111111111111110101110001, 24'b111111111111111111111111, 24'b000000000000000100110000, 24'b111111111111111111111111, 24'b000000000000000010000100, 24'b111111111111111111101100, 24'b000000000000000100010100, 24'b000000000000000000000000, 24'b000000000000000101010100, 24'b111111111111100111101101, 24'b111111111111111111111111}, 
{24'b000000000000010011110111, 24'b111111111111111111011011, 24'b000000000000001001100110, 24'b111111111111101100011101, 24'b111111111111110011101001, 24'b111111111111111111111111, 24'b111111111111111111111111, 24'b000000000000000001110000, 24'b000000000000000000001001, 24'b111111111111110111111100, 24'b000000000000000000000000, 24'b000000000000000000001000, 24'b000000000000000000000000, 24'b000000000000000000000001, 24'b111111111111110111101111, 24'b000000000000001001001000, 24'b111111111111111111111001, 24'b111111111111111110000001, 24'b000000000000000000000000, 24'b000000000000000111101011, 24'b111111111111110011001001, 24'b000000000000000111011011, 24'b000000000000001000111101, 24'b000000000000001000010000, 24'b111111111111111111111111, 24'b000000000000100011010010, 24'b111111111111110110001100, 24'b000000000000010111010000, 24'b111111111111111100101100, 24'b111111111111101000111010, 24'b111111111111110100111001, 24'b000000000000001000111011}, 
{24'b111111111111011101001111, 24'b111111111111111110010010, 24'b111111111111110110001001, 24'b111111111111111111111111, 24'b000000000000010000101100, 24'b111111111111110100100100, 24'b111111111111111100001010, 24'b000000000000001111001111, 24'b000000000000000110000011, 24'b111111111111110000110001, 24'b000000000000000000000000, 24'b111111111111111110001100, 24'b111111111111111111010111, 24'b000000000000001000110011, 24'b111111111111110000010001, 24'b111111111111111111010010, 24'b000000000000000000000000, 24'b111111111111111111111101, 24'b111111111111111110111110, 24'b000000000000000000000000, 24'b111111111111110011110101, 24'b111111111111111111111111, 24'b000000000000000000000000, 24'b111111111111101010111111, 24'b000000000000000100011111, 24'b000000000000100111101010, 24'b000000000000010110001000, 24'b111111111111111101101101, 24'b111111111111110101101110, 24'b111111111111100011010010, 24'b000000000000000000000001, 24'b111111111111111100111000}, 
{24'b000000000000000001010111, 24'b000000000000001101101011, 24'b000000000000000001010111, 24'b111111111111110110010101, 24'b000000000000000000010010, 24'b111111111111111110010111, 24'b000000000000000000000000, 24'b000000000000001101010101, 24'b000000000000001101110000, 24'b111111111111110111011100, 24'b000000000000001000111111, 24'b000000000000000001100010, 24'b111111111111111111111111, 24'b111111111111111111000101, 24'b111111111111110101110101, 24'b000000000000010000001100, 24'b111111111111111101010010, 24'b111111111111101011010100, 24'b000000000000000111010100, 24'b111111111111111111111111, 24'b111111111111111111111111, 24'b000000000000000111011110, 24'b111111111111111011001111, 24'b111111111111111111101100, 24'b111111111111111100101100, 24'b000000000000000101101001, 24'b111111111111110111000001, 24'b000000000000001000100101, 24'b111111111111101000101110, 24'b000000000000000101001001, 24'b111111111111111111111110, 24'b000000000000001010000001}, 
{24'b111111111111111101010000, 24'b000000000000000000000010, 24'b000000000000000101101100, 24'b000000000000000000000000, 24'b111111111111111100000110, 24'b111111111111111111110100, 24'b000000000000000110100100, 24'b111111111111111111111111, 24'b000000000000000000000000, 24'b000000000000000000010100, 24'b000000000000000000000000, 24'b000000000000000001010001, 24'b111111111111111001001100, 24'b000000000000000000101010, 24'b000000000000000111000101, 24'b000000000000000010111111, 24'b000000000000000110110000, 24'b111111111111111111111101, 24'b111111111111111111111010, 24'b000000000000001000001100, 24'b000000000000001111110101, 24'b111111111111111001101111, 24'b000000000000000000000000, 24'b111111111111111111110111, 24'b000000000000000000101110, 24'b111111111111100010011111, 24'b111111111111111111111100, 24'b111111111111111011011110, 24'b111111111111111111111111, 24'b000000000000100100001000, 24'b000000000000000000000001, 24'b111111111111110010110100}, 
{24'b111111111111111110010010, 24'b111111111111111000010111, 24'b111111111111111111011011, 24'b000000000000000000011100, 24'b000000000000000101110011, 24'b111111111111111111111111, 24'b000000000000000000000000, 24'b111111111111111110100001, 24'b000000000000000100100001, 24'b111111111111111111011110, 24'b000000000000000000000000, 24'b000000000000000010000001, 24'b000000000000010010111000, 24'b111111111111111001011110, 24'b000000000000000000110011, 24'b111111111111001001101101, 24'b111111111111111111010010, 24'b111111111111111100001000, 24'b000000000000000000100000, 24'b111111111111111100110011, 24'b000000000000000101111000, 24'b111111111111110001101010, 24'b000000000000000111010011, 24'b000000000000000110101111, 24'b111111111111111111001010, 24'b111111111111010010011111, 24'b111111111111110001010111, 24'b111111111111111110100110, 24'b111111111111111110110100, 24'b000000000000011000111111, 24'b111111111111111111101000, 24'b000000000000001001110111}, 
{24'b000000000000000011000000, 24'b000000000000000000000000, 24'b000000000000001011001001, 24'b111111111111111000101111, 24'b111111111111111011100110, 24'b000000000000001111001110, 24'b111111111111110101110001, 24'b000000000000000011101011, 24'b111111111111101100001100, 24'b000000000000000000100011, 24'b000000000000000001000100, 24'b111111111111111010101000, 24'b000000000000000000000010, 24'b000000000000000000000000, 24'b111111111111110011111110, 24'b000000000000011011101011, 24'b111111111111110000001101, 24'b111111111111111111001111, 24'b000000000000000111100110, 24'b111111111111111111111111, 24'b000000000000000100011011, 24'b111111111111100001010101, 24'b000000000000010100000010, 24'b111111111111111111111111, 24'b111111111111111000000100, 24'b000000000000011111000001, 24'b000000000000001001010110, 24'b111111111111110101111001, 24'b111111111111110111011001, 24'b111111111111011101100111, 24'b111111111111111111010110, 24'b000000000000000001000001}, 
{24'b111111111111111111111111, 24'b000000000000000000011010, 24'b111111111111111101110001, 24'b111111111111101110110110, 24'b111111111111111111111110, 24'b111111111111100110111000, 24'b000000000000000000000001, 24'b000000000000010011011011, 24'b000000000000001111101000, 24'b000000000000000001001101, 24'b000000000000000000000000, 24'b111111111111111000111100, 24'b000000000000010101010000, 24'b111111111111111111111111, 24'b111111111111111111111110, 24'b111111111111111111111110, 24'b000000000000011011110001, 24'b000000000000000000000110, 24'b111111111111111101011101, 24'b111111111111111100101110, 24'b111111111111101011011001, 24'b000000000000001000011011, 24'b000000000000000000000000, 24'b000000000000000000000000, 24'b000000000000000010000001, 24'b111111111111111011011100, 24'b111111111111100010100001, 24'b000000000000010001101010, 24'b111111111111100011100111, 24'b000000000000000011010001, 24'b111111111111111010111100, 24'b000000000000000000000000}, 
{24'b000000000000000011111011, 24'b000000000000001011111011, 24'b000000000000000000100111, 24'b111111111111111111110011, 24'b111111111111100010100110, 24'b000000000000000000000011, 24'b111111111111111111111111, 24'b000000000000001111100000, 24'b000000000000010001101110, 24'b111111111111111111111111, 24'b111111111111111111111111, 24'b111111111111111111111010, 24'b000000000000000000000000, 24'b000000000000000000001000, 24'b000000000000000000000000, 24'b000000000000000000000000, 24'b000000000000000000000001, 24'b111111111111111111111101, 24'b000000000000001010111000, 24'b111111111111111001011010, 24'b111111111111100100010110, 24'b111111111111111101111000, 24'b111111111111111001101011, 24'b111111111111111001111111, 24'b111111111111111011100100, 24'b111111111111111111111100, 24'b111111111111111011111110, 24'b111111111111111110100110, 24'b111111111111111111010101, 24'b000000000000001001000011, 24'b111111111111111111111110, 24'b000000000000011101101010}
};

localparam logic signed [23:0] bias [32] = '{
24'b000000000001011110010110,  // 1.474280834197998
24'b000000000000101100010000,  // 0.6914801001548767
24'b000000000001011100001100,  // 1.4406442642211914
24'b000000000001011010000111,  // 1.408045768737793
24'b000000000000111111001000,  // 0.9864811301231384
24'b000000000000110111010001,  // 0.8636202812194824
24'b111111111111011000100111,  // -0.6153604388237
24'b000000000000011110111110,  // 0.4839226007461548
24'b000000000000011111000111,  // 0.4862793982028961
24'b000000000000010111110010,  // 0.37162142992019653
24'b000000000000011101011011,  // 0.45989668369293213
24'b000000000001010011001100,  // 1.2998151779174805
24'b111111111110111110111100,  // -1.016528844833374
24'b111111111111101001011100,  // -0.35249894857406616
24'b000000000000011100100010,  // 0.44582197070121765
24'b111111111111111000110101,  // -0.1119980737566948
24'b111111111111111011101100,  // -0.06717441976070404
24'b000000000000000000010011,  // 0.00487547367811203
24'b000000000000001100011101,  // 0.1946917623281479
24'b111111111111001110000110,  // -0.7796769738197327
24'b000000000000101110101000,  // 0.7287401556968689
24'b000000000001101101110000,  // 1.714877724647522
24'b111111111110011001110010,  // -1.5971007347106934
24'b000000000000000100101110,  // 0.07393483817577362
24'b000000000000010100101001,  // 0.3225609362125397
24'b000000000000110110000110,  // 0.8453295230865479
24'b000000000000111001100000,  // 0.898597240447998
24'b000000000000010000010011,  // 0.2548799514770508
24'b000000000000111110010011,  // 0.9735668301582336
24'b000000000001001000000100,  // 1.1261906623840332
24'b000000000000011100101001,  // 0.44768181443214417
24'b111111111101101000011110   // -2.3676068782806396
};
endpackage