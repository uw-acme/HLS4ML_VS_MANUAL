// Package with weights and biases for pre-sigmoid dense latency layer
`ifndef DENSE_LAYER_1_PKG
    `define DENSE_LAYER_1_PKG dense_1_16_10
`endif

`ifndef DENSE_LAYER_2_PKG
    `define DENSE_LAYER_2_PKG dense_2_16_10
`endif

`ifndef DENSE_LAYER_3_PKG
    `define DENSE_LAYER_3_PKG dense_3_16_10
`endif

`ifndef DENSE_LAYER_4_PKG
    `define DENSE_LAYER_4_PKG dense_4_16_10
`endif