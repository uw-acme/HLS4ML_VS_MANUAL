// Width: 19
// NFRAC: 9
package dense_4_19_9;

localparam logic signed [18:0] weights [32][5] = '{ 
{19'b1111111111111111001, 19'b0000000000010100001, 19'b1111111111101100111, 19'b0000000000000100001, 19'b1111111111111001001}, 
{19'b1111111111011100010, 19'b1111111111111100011, 19'b0000000000011101011, 19'b1111111111111111001, 19'b0000000000000001000}, 
{19'b0000000000010111110, 19'b0000000000001101100, 19'b1111111111111110001, 19'b1111111111100110000, 19'b1111111111110010100}, 
{19'b1111111111100111111, 19'b1111111111101000001, 19'b1111111111111000110, 19'b0000000000010011101, 19'b0000000000001111000}, 
{19'b0000000000000111110, 19'b0000000000001000001, 19'b0000000000001010000, 19'b1111111111111110110, 19'b1111111110111111001}, 
{19'b0000000000010100111, 19'b1111111111100110110, 19'b0000000000001011100, 19'b1111111111110101101, 19'b1111111111110101000}, 
{19'b1111111111100110010, 19'b0000000000000010010, 19'b1111111111111111111, 19'b0000000000001011001, 19'b0000000000000100011}, 
{19'b1111111111111111111, 19'b0000000000010010001, 19'b1111111111100110111, 19'b0000000000001010011, 19'b0000000000001000101}, 
{19'b0000000000001010011, 19'b1111111111110101001, 19'b0000000000000000000, 19'b1111111111100010011, 19'b1111111111110000000}, 
{19'b1111111111111111111, 19'b1111111111101110111, 19'b0000000000001011011, 19'b0000000000011011100, 19'b0000000000000000000}, 
{19'b1111111111110111101, 19'b1111111111110110101, 19'b0000000000000000000, 19'b0000000000100101001, 19'b1111111111101110110}, 
{19'b0000000000001010110, 19'b0000000000001110101, 19'b1111111111101010001, 19'b1111111111111110001, 19'b0000000000000111110}, 
{19'b0000000000000000000, 19'b0000000000001010101, 19'b0000000000000000100, 19'b1111111111110010101, 19'b1111111111011000001}, 
{19'b0000000000001011010, 19'b0000000000000100000, 19'b0000000000011010110, 19'b1111111111111011100, 19'b1111111111100100100}, 
{19'b0000000000000101110, 19'b1111111111111100111, 19'b1111111111101000111, 19'b1111111111111101111, 19'b0000000000100010010}, 
{19'b1111111111100001101, 19'b1111111111110000010, 19'b1111111111110001110, 19'b0000000000011001100, 19'b0000000000000010000}, 
{19'b0000000000010110001, 19'b1111111111110101000, 19'b1111111111110111010, 19'b1111111111110001100, 19'b1111111111111100001}, 
{19'b0000000000001100011, 19'b1111111111111101011, 19'b1111111111100101100, 19'b1111111111111110000, 19'b0000000000000100100}, 
{19'b0000000000010000100, 19'b0000000000000010101, 19'b1111111111110010000, 19'b0000000000000000000, 19'b1111111111100111111}, 
{19'b0000000000001110110, 19'b1111111111111010011, 19'b1111111111110010011, 19'b0000000000001101010, 19'b0000000000000110000}, 
{19'b0000000000000100010, 19'b1111111111111110000, 19'b0000000000010011000, 19'b1111111111100100011, 19'b1111111111111110101}, 
{19'b0000000000000000000, 19'b0000000000000111100, 19'b0000000000011111001, 19'b1111111111011110110, 19'b1111111111011000011}, 
{19'b1111111111111001101, 19'b0000000000000111000, 19'b0000000000001011010, 19'b1111111111101001001, 19'b0000000000100001011}, 
{19'b1111111111111111111, 19'b0000000000001010100, 19'b0000000000010010000, 19'b0000000000000010011, 19'b1111111111011011011}, 
{19'b1111111111110101001, 19'b0000000000010111010, 19'b1111111111110001101, 19'b0000000000000000010, 19'b0000000000011000110}, 
{19'b0000000000000001101, 19'b0000000000010001000, 19'b0000000000000001111, 19'b1111111111010000001, 19'b0000000000100011000}, 
{19'b1111111111100010100, 19'b1111111111110000011, 19'b0000000000001101101, 19'b0000000000001111101, 19'b0000000000001100111}, 
{19'b0000000000000000010, 19'b0000000000001111011, 19'b1111111111111101101, 19'b1111111111110110010, 19'b0000000000000010000}, 
{19'b1111111111111001010, 19'b0000000000001111110, 19'b1111111111011111110, 19'b0000000000001000111, 19'b1111111111110101110}, 
{19'b1111111111111110110, 19'b0000000000001001000, 19'b1111111111110101001, 19'b1111111111100110010, 19'b0000000000100101111}, 
{19'b0000000000011100101, 19'b0000000000000100011, 19'b0000000000010100110, 19'b1111111111011010010, 19'b1111111111101011110}, 
{19'b1111111111111100001, 19'b1111111111100111010, 19'b0000000000010111011, 19'b0000000000000100100, 19'b0000000000001000001}
};

localparam logic signed [18:0] bias [5] = '{
19'b1111111111111100000,  // -0.06223141402006149
19'b1111111111111011111,  // -0.06270556896924973
19'b1111111111111011100,  // -0.07014333456754684
19'b0000000000000101010,  // 0.0820775106549263
19'b0000000000001101110   // 0.2155742198228836
};
endpackage