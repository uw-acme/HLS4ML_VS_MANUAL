// Width: 6
// NFRAC: 3
package dense_2_6_3;

localparam logic signed [5:0] weights [64][32] = '{ 
{6'b000010, 6'b000000, 6'b111110, 6'b111111, 6'b000010, 6'b000000, 6'b111110, 6'b111111, 6'b111101, 6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b111110, 6'b111111, 6'b111101, 6'b000000, 6'b111111, 6'b111110, 6'b111110, 6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b000011, 6'b000001, 6'b111111, 6'b000000, 6'b111100, 6'b000000}, 
{6'b111111, 6'b111110, 6'b111110, 6'b111111, 6'b111111, 6'b000000, 6'b111110, 6'b000000, 6'b000000, 6'b111111, 6'b000001, 6'b111111, 6'b111111, 6'b111110, 6'b000000, 6'b111111, 6'b000000, 6'b111110, 6'b000001, 6'b000001, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b000010, 6'b000001, 6'b000000, 6'b000000, 6'b111100, 6'b000000, 6'b000000}, 
{6'b000000, 6'b111111, 6'b111110, 6'b111111, 6'b111111, 6'b111111, 6'b111110, 6'b000000, 6'b111110, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b000001, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b000001, 6'b000001, 6'b000000, 6'b111111, 6'b111110, 6'b111111, 6'b000000}, 
{6'b000001, 6'b000000, 6'b000000, 6'b111111, 6'b111011, 6'b000000, 6'b000000, 6'b000001, 6'b000001, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b000001, 6'b000000, 6'b111111, 6'b111111, 6'b111110, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b111110, 6'b000010}, 
{6'b111010, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b111110, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b000001, 6'b000000, 6'b000010, 6'b111111, 6'b000001, 6'b111100, 6'b000000, 6'b111111, 6'b000001, 6'b000010, 6'b000000, 6'b000000, 6'b000001, 6'b000001, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b000001}, 
{6'b000000, 6'b111111, 6'b000001, 6'b111010, 6'b110100, 6'b111101, 6'b000010, 6'b111011, 6'b111111, 6'b111010, 6'b111011, 6'b111101, 6'b000010, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b111110, 6'b111111, 6'b111100, 6'b000000, 6'b000001, 6'b111111, 6'b000000, 6'b000010, 6'b000000, 6'b111111, 6'b111111, 6'b000001, 6'b111111, 6'b000001}, 
{6'b111111, 6'b111110, 6'b111110, 6'b111111, 6'b111101, 6'b000000, 6'b111110, 6'b111110, 6'b111100, 6'b000000, 6'b111111, 6'b111110, 6'b000000, 6'b111111, 6'b111111, 6'b111011, 6'b111111, 6'b000000, 6'b000001, 6'b111110, 6'b111110, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b111010, 6'b111101, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b111111}, 
{6'b111110, 6'b111111, 6'b111111, 6'b111110, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b000001, 6'b000000, 6'b000000, 6'b111111, 6'b000001, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b111110, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b111111}, 
{6'b111100, 6'b111111, 6'b111100, 6'b000000, 6'b000011, 6'b111111, 6'b111111, 6'b000001, 6'b111100, 6'b111111, 6'b000000, 6'b111110, 6'b111111, 6'b000000, 6'b111110, 6'b000110, 6'b111111, 6'b000000, 6'b000001, 6'b000001, 6'b000000, 6'b111101, 6'b000000, 6'b000011, 6'b111110, 6'b000101, 6'b111110, 6'b111110, 6'b111100, 6'b111100, 6'b000000, 6'b000000}, 
{6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b000010, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b111110, 6'b000000, 6'b000001, 6'b111111, 6'b000000, 6'b000000, 6'b000000}, 
{6'b000000, 6'b000000, 6'b111111, 6'b111101, 6'b111001, 6'b000001, 6'b000000, 6'b111001, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b111100, 6'b111111, 6'b000001, 6'b000001, 6'b000001, 6'b111100, 6'b111101, 6'b000000, 6'b111111, 6'b111111, 6'b000010, 6'b111111, 6'b111111, 6'b111111, 6'b000001, 6'b111111, 6'b000000}, 
{6'b111110, 6'b111100, 6'b000000, 6'b111111, 6'b000010, 6'b111101, 6'b111110, 6'b000000, 6'b111111, 6'b000001, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b111101, 6'b000001, 6'b000000, 6'b000010, 6'b000000, 6'b000000, 6'b111111, 6'b000001, 6'b111111, 6'b111101, 6'b111111, 6'b000001, 6'b111111, 6'b000000, 6'b111111, 6'b000001, 6'b000010}, 
{6'b000000, 6'b000000, 6'b000001, 6'b000000, 6'b111111, 6'b000001, 6'b000000, 6'b111111, 6'b000000, 6'b111110, 6'b111111, 6'b111110, 6'b111111, 6'b000000, 6'b111111, 6'b000110, 6'b000000, 6'b111111, 6'b111110, 6'b111111, 6'b000001, 6'b000001, 6'b000000, 6'b111111, 6'b000001, 6'b000010, 6'b000011, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b111111}, 
{6'b111110, 6'b000000, 6'b000000, 6'b111110, 6'b111101, 6'b000011, 6'b000000, 6'b000000, 6'b111110, 6'b111111, 6'b000001, 6'b000000, 6'b000000, 6'b111111, 6'b000010, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b000101, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b000001}, 
{6'b000000, 6'b000000, 6'b000010, 6'b111111, 6'b000000, 6'b000010, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b000011, 6'b111111, 6'b000000, 6'b000001, 6'b000000, 6'b000000, 6'b111101, 6'b111110, 6'b111111, 6'b111111, 6'b111110, 6'b111111, 6'b111111, 6'b111110, 6'b111110, 6'b000000, 6'b000000, 6'b111100, 6'b000000}, 
{6'b111101, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b000001, 6'b111111, 6'b000010, 6'b111101, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b000001, 6'b111111, 6'b111101, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b111110, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b111110}, 
{6'b111101, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000001, 6'b000000, 6'b111111, 6'b000000, 6'b000011, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b000001, 6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b111110, 6'b000001, 6'b111111, 6'b000000, 6'b111110}, 
{6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b000111, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b000001, 6'b000000, 6'b111110, 6'b111111, 6'b111111, 6'b000010, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b000000}, 
{6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b000010, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b111110, 6'b111110, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b111110, 6'b000000, 6'b111110, 6'b000000, 6'b000000, 6'b111110, 6'b000000, 6'b000000, 6'b111111}, 
{6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b000001, 6'b111111, 6'b111111, 6'b000000, 6'b111100, 6'b000000, 6'b111111, 6'b111111, 6'b000010, 6'b000001, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b111110, 6'b111111, 6'b000001, 6'b000000, 6'b111110, 6'b000000, 6'b111111, 6'b111111, 6'b000001, 6'b000000, 6'b111110}, 
{6'b000101, 6'b000010, 6'b111110, 6'b000000, 6'b111101, 6'b000000, 6'b000001, 6'b000000, 6'b000001, 6'b111111, 6'b111110, 6'b111111, 6'b000001, 6'b000000, 6'b111111, 6'b000001, 6'b000100, 6'b111110, 6'b111101, 6'b000000, 6'b111111, 6'b111110, 6'b111111, 6'b111111, 6'b000000, 6'b111101, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b000000}, 
{6'b111111, 6'b111110, 6'b111111, 6'b111110, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b111110, 6'b000000, 6'b000000, 6'b111111, 6'b000011, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b000010, 6'b111100, 6'b111111, 6'b111111, 6'b111111, 6'b000001, 6'b111111, 6'b000000, 6'b000011, 6'b111011, 6'b111101, 6'b000000}, 
{6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b111010, 6'b111011, 6'b000000, 6'b111111, 6'b111101, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b111110, 6'b000010, 6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b000001, 6'b111011, 6'b000001, 6'b111111, 6'b111111, 6'b000001, 6'b111111, 6'b000001}, 
{6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b111101, 6'b000000, 6'b000000, 6'b000100, 6'b111111, 6'b000000, 6'b000000, 6'b000010, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b111101, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b000001, 6'b000000, 6'b000001, 6'b111100, 6'b000000, 6'b000011, 6'b000000}, 
{6'b111101, 6'b000001, 6'b111101, 6'b000000, 6'b111111, 6'b000000, 6'b000011, 6'b111110, 6'b111101, 6'b000001, 6'b111110, 6'b111111, 6'b111111, 6'b000010, 6'b111111, 6'b111101, 6'b111111, 6'b000011, 6'b111100, 6'b111111, 6'b000010, 6'b111101, 6'b000000, 6'b111111, 6'b000010, 6'b111011, 6'b111101, 6'b111110, 6'b111111, 6'b000000, 6'b000000, 6'b000001}, 
{6'b111111, 6'b000000, 6'b111111, 6'b000001, 6'b111111, 6'b000001, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b000100, 6'b000000, 6'b000001, 6'b000000, 6'b111110, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b111110, 6'b111111, 6'b000010, 6'b000010, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b111111}, 
{6'b111111, 6'b000000, 6'b000010, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b111001, 6'b000001, 6'b000000, 6'b000000, 6'b111101, 6'b000000, 6'b111110, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b000010, 6'b000011, 6'b111110, 6'b111110, 6'b000001, 6'b111101, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b000001}, 
{6'b111111, 6'b111111, 6'b111110, 6'b111110, 6'b111111, 6'b111110, 6'b000000, 6'b000000, 6'b111110, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b000001, 6'b000001, 6'b111110, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b111101, 6'b111111, 6'b000001}, 
{6'b111111, 6'b111111, 6'b000000, 6'b000010, 6'b000000, 6'b000000, 6'b000000, 6'b111110, 6'b111110, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000001, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b000001, 6'b000000, 6'b111111, 6'b111110, 6'b111111, 6'b111101, 6'b000000, 6'b000000, 6'b000000}, 
{6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b111110, 6'b111110, 6'b000000, 6'b000000, 6'b111110, 6'b000001, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b111110, 6'b000000, 6'b111110, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000010, 6'b000000, 6'b000000, 6'b000000}, 
{6'b111111, 6'b000010, 6'b111111, 6'b111111, 6'b111110, 6'b111111, 6'b000011, 6'b111010, 6'b111101, 6'b111110, 6'b111110, 6'b111101, 6'b111111, 6'b000011, 6'b111111, 6'b000000, 6'b111110, 6'b000011, 6'b111100, 6'b000000, 6'b111111, 6'b111101, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b111110, 6'b111111, 6'b000001, 6'b000000, 6'b111111, 6'b000000}, 
{6'b000010, 6'b111111, 6'b000001, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b000001, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b111101, 6'b111111, 6'b000000, 6'b111111, 6'b111110, 6'b111111, 6'b111111, 6'b000100, 6'b111101, 6'b111111}, 
{6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b000001, 6'b111110, 6'b111111, 6'b111110, 6'b000000, 6'b000001, 6'b111110, 6'b111101, 6'b000000, 6'b111010, 6'b111111, 6'b111111, 6'b111110, 6'b111111, 6'b000001, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b111001, 6'b111011, 6'b111101, 6'b000000, 6'b000001, 6'b111111, 6'b000001}, 
{6'b111111, 6'b111110, 6'b000001, 6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b000100, 6'b111110, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b000001, 6'b111110, 6'b111111, 6'b000001, 6'b111111, 6'b000000, 6'b000100, 6'b000010, 6'b000000, 6'b000000, 6'b111100, 6'b111111, 6'b111111}, 
{6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b000001, 6'b111100, 6'b000000, 6'b111111, 6'b000001, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b000010, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b111101, 6'b000000, 6'b000001, 6'b111111, 6'b000000, 6'b111111, 6'b000000}, 
{6'b111110, 6'b000000, 6'b111100, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b111110, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b000010, 6'b111111, 6'b000000, 6'b111111, 6'b000010, 6'b000001, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b000000}, 
{6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b111100, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b111110, 6'b111111, 6'b000000, 6'b111110, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b111101, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b000001, 6'b111111, 6'b000000, 6'b000011, 6'b000010, 6'b000000, 6'b000000, 6'b111110, 6'b000000, 6'b111111}, 
{6'b000000, 6'b000000, 6'b000010, 6'b111110, 6'b000001, 6'b000000, 6'b000000, 6'b000001, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b111011, 6'b111111, 6'b000000, 6'b111111, 6'b111011, 6'b111110, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b111111}, 
{6'b000000, 6'b111111, 6'b111111, 6'b111110, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b000001, 6'b111111, 6'b000000, 6'b111101, 6'b111111, 6'b000001, 6'b111111, 6'b111101, 6'b000000, 6'b111111, 6'b000010, 6'b111111, 6'b111100, 6'b111111, 6'b000010, 6'b111111, 6'b111111, 6'b000001, 6'b111111, 6'b000000, 6'b000000, 6'b111110, 6'b000000, 6'b000000}, 
{6'b111110, 6'b000000, 6'b000000, 6'b111111, 6'b000011, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b000001, 6'b111111, 6'b000001, 6'b000000, 6'b111111, 6'b111101, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b111110, 6'b111101, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b000000}, 
{6'b111100, 6'b111110, 6'b111110, 6'b000000, 6'b000100, 6'b111110, 6'b000000, 6'b111111, 6'b111100, 6'b000001, 6'b111111, 6'b000100, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b000011, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b111100, 6'b111110, 6'b111111, 6'b111111, 6'b111111}, 
{6'b000001, 6'b111001, 6'b111010, 6'b111110, 6'b000101, 6'b111111, 6'b111101, 6'b000010, 6'b000000, 6'b000000, 6'b000001, 6'b111101, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b111000, 6'b000001, 6'b000010, 6'b000010, 6'b000000, 6'b000000, 6'b111100, 6'b111010, 6'b111111, 6'b111101, 6'b111100, 6'b111110, 6'b111000, 6'b000011, 6'b000011}, 
{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000010, 6'b111110, 6'b000000, 6'b000000, 6'b111101, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b000001, 6'b000000, 6'b000000, 6'b000000, 6'b000010, 6'b111110, 6'b000000, 6'b111110, 6'b111111, 6'b000010, 6'b000000, 6'b111111, 6'b111011, 6'b111111, 6'b111110, 6'b111111, 6'b000000, 6'b000001, 6'b000000}, 
{6'b111111, 6'b000001, 6'b111101, 6'b000000, 6'b000001, 6'b111111, 6'b111111, 6'b000001, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b000011, 6'b000000, 6'b111101, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b000010, 6'b111111}, 
{6'b111111, 6'b000000, 6'b111111, 6'b111110, 6'b111001, 6'b000000, 6'b000000, 6'b111111, 6'b111011, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b111101, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b000010, 6'b111111, 6'b111101, 6'b000000, 6'b111101, 6'b111111, 6'b111110, 6'b111111, 6'b111111, 6'b111111, 6'b111100, 6'b111111, 6'b000001}, 
{6'b000000, 6'b000001, 6'b111111, 6'b000001, 6'b111110, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b111101, 6'b111111, 6'b000001, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b000001, 6'b111101, 6'b000010, 6'b000000, 6'b000000, 6'b000001, 6'b000000, 6'b111111, 6'b111100, 6'b111111, 6'b111110, 6'b000001}, 
{6'b000000, 6'b000000, 6'b111101, 6'b111111, 6'b000001, 6'b111110, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b111110, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b111110, 6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b000010, 6'b111111, 6'b000000, 6'b111101, 6'b111101, 6'b000001, 6'b111111, 6'b111111, 6'b000000, 6'b000010}, 
{6'b111101, 6'b111111, 6'b111110, 6'b000000, 6'b111101, 6'b000000, 6'b111111, 6'b111111, 6'b111011, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b111110, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b000010, 6'b111111, 6'b000001, 6'b000000, 6'b111110, 6'b000001, 6'b111111, 6'b000000, 6'b111111, 6'b000100}, 
{6'b111101, 6'b000000, 6'b000000, 6'b111111, 6'b000001, 6'b111101, 6'b111111, 6'b000010, 6'b000001, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b000001, 6'b000000, 6'b000000, 6'b000000, 6'b000010, 6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b000000}, 
{6'b111111, 6'b000000, 6'b111110, 6'b111111, 6'b000010, 6'b111111, 6'b111111, 6'b000001, 6'b111111, 6'b000010, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b111101, 6'b000010, 6'b000001, 6'b000101, 6'b000001, 6'b000001, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b111100, 6'b111111, 6'b111111, 6'b111111}, 
{6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b111110, 6'b000000, 6'b000001, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b000001, 6'b111111, 6'b111111, 6'b111101, 6'b000000, 6'b111110, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b000001, 6'b111111, 6'b111111, 6'b111100, 6'b000000}, 
{6'b000011, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b000001, 6'b000000, 6'b000100, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b111100, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b111101, 6'b111111, 6'b000001, 6'b111111, 6'b000010, 6'b111111, 6'b111110}, 
{6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b111101, 6'b111111, 6'b000000, 6'b111111, 6'b000001, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b000010, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b000001, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b000000}, 
{6'b111101, 6'b000001, 6'b000000, 6'b111111, 6'b111100, 6'b111111, 6'b000000, 6'b111100, 6'b000100, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b111100, 6'b000000, 6'b000001, 6'b000000, 6'b000000, 6'b111010, 6'b111101, 6'b111110, 6'b000000, 6'b111111, 6'b000010, 6'b111110}, 
{6'b111111, 6'b111110, 6'b111111, 6'b111100, 6'b111101, 6'b000010, 6'b000010, 6'b111110, 6'b000000, 6'b111111, 6'b111111, 6'b111101, 6'b000000, 6'b111101, 6'b000001, 6'b111111, 6'b000010, 6'b111111, 6'b111111, 6'b111110, 6'b111111, 6'b111111, 6'b111101, 6'b000000, 6'b111111, 6'b111111, 6'b111110, 6'b000010, 6'b000010, 6'b111111, 6'b111010, 6'b000001}, 
{6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b111110, 6'b111111, 6'b000000, 6'b000001, 6'b000000, 6'b000001, 6'b111111, 6'b111110, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b111100, 6'b111111}, 
{6'b000010, 6'b111111, 6'b000001, 6'b111101, 6'b111110, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b111110, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b111110, 6'b000001, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b111110, 6'b000000, 6'b000001, 6'b000001, 6'b111111, 6'b000100, 6'b111110, 6'b000010, 6'b111111, 6'b111101, 6'b111110, 6'b000001}, 
{6'b111011, 6'b111111, 6'b111110, 6'b111111, 6'b000010, 6'b111110, 6'b111111, 6'b000001, 6'b000000, 6'b111110, 6'b000000, 6'b111111, 6'b111111, 6'b000001, 6'b111110, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b111110, 6'b111111, 6'b000000, 6'b111101, 6'b000000, 6'b000100, 6'b000010, 6'b111111, 6'b111110, 6'b111100, 6'b000000, 6'b111111}, 
{6'b000000, 6'b000001, 6'b000000, 6'b111110, 6'b000000, 6'b111111, 6'b000000, 6'b000001, 6'b000001, 6'b111110, 6'b000001, 6'b000000, 6'b111111, 6'b111111, 6'b111110, 6'b000010, 6'b111111, 6'b111101, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b111110, 6'b000001, 6'b111101, 6'b000000, 6'b111111, 6'b000001}, 
{6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b111111, 6'b000001, 6'b000001, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b111100, 6'b111111, 6'b111111, 6'b111111, 6'b000100, 6'b000000, 6'b111110}, 
{6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b000010, 6'b111111, 6'b000000, 6'b111001, 6'b111111, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b111110, 6'b000000, 6'b000000, 6'b111111, 6'b111010, 6'b111110, 6'b111111, 6'b111111, 6'b000011, 6'b111111, 6'b000001}, 
{6'b000000, 6'b000000, 6'b000001, 6'b111111, 6'b111111, 6'b000001, 6'b111110, 6'b000000, 6'b111101, 6'b000000, 6'b000000, 6'b111111, 6'b000000, 6'b000000, 6'b111110, 6'b000011, 6'b111110, 6'b111111, 6'b000000, 6'b111111, 6'b000000, 6'b111100, 6'b000010, 6'b111111, 6'b111111, 6'b000011, 6'b000001, 6'b111110, 6'b111110, 6'b111011, 6'b111111, 6'b000000}, 
{6'b111111, 6'b000000, 6'b111111, 6'b111101, 6'b111111, 6'b111100, 6'b000000, 6'b000010, 6'b000001, 6'b000000, 6'b000000, 6'b111111, 6'b000010, 6'b111111, 6'b111111, 6'b111111, 6'b000011, 6'b000000, 6'b111111, 6'b111111, 6'b111101, 6'b000001, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b111100, 6'b000010, 6'b111100, 6'b000000, 6'b111111, 6'b000000}, 
{6'b000000, 6'b000001, 6'b000000, 6'b111111, 6'b111100, 6'b000000, 6'b111111, 6'b000001, 6'b000010, 6'b111111, 6'b111111, 6'b111111, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b111111, 6'b000001, 6'b111111, 6'b111100, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b111111, 6'b000001, 6'b111111, 6'b000011}
};

localparam logic signed [5:0] bias [32] = '{
6'b001011,  // 1.474280834197998
6'b000101,  // 0.6914801001548767
6'b001011,  // 1.4406442642211914
6'b001011,  // 1.408045768737793
6'b000111,  // 0.9864811301231384
6'b000110,  // 0.8636202812194824
6'b111011,  // -0.6153604388237
6'b000011,  // 0.4839226007461548
6'b000011,  // 0.4862793982028961
6'b000010,  // 0.37162142992019653
6'b000011,  // 0.45989668369293213
6'b001010,  // 1.2998151779174805
6'b110111,  // -1.016528844833374
6'b111101,  // -0.35249894857406616
6'b000011,  // 0.44582197070121765
6'b111111,  // -0.1119980737566948
6'b111111,  // -0.06717441976070404
6'b000000,  // 0.00487547367811203
6'b000001,  // 0.1946917623281479
6'b111001,  // -0.7796769738197327
6'b000101,  // 0.7287401556968689
6'b001101,  // 1.714877724647522
6'b110011,  // -1.5971007347106934
6'b000000,  // 0.07393483817577362
6'b000010,  // 0.3225609362125397
6'b000110,  // 0.8453295230865479
6'b000111,  // 0.898597240447998
6'b000010,  // 0.2548799514770508
6'b000111,  // 0.9735668301582336
6'b001001,  // 1.1261906623840332
6'b000011,  // 0.44768181443214417
6'b101101   // -2.3676068782806396
};
endpackage