// Width: 21
// NFRAC: 10
package dense_4_21_10;

localparam logic signed [20:0] weights [32][5] = '{ 
{21'b111111111111111110011, 21'b000000000000101000011, 21'b111111111111011001110, 21'b000000000000001000011, 21'b111111111111110010011}, 
{21'b111111111110111000100, 21'b111111111111111000111, 21'b000000000000111010111, 21'b111111111111111110011, 21'b000000000000000010001}, 
{21'b000000000000101111100, 21'b000000000000011011000, 21'b111111111111111100011, 21'b111111111111001100000, 21'b111111111111100101000}, 
{21'b111111111111001111111, 21'b111111111111010000010, 21'b111111111111110001101, 21'b000000000000100111011, 21'b000000000000011110000}, 
{21'b000000000000001111101, 21'b000000000000010000011, 21'b000000000000010100000, 21'b111111111111111101101, 21'b111111111101111110010}, 
{21'b000000000000101001110, 21'b111111111111001101100, 21'b000000000000010111001, 21'b111111111111101011010, 21'b111111111111101010001}, 
{21'b111111111111001100101, 21'b000000000000000100100, 21'b111111111111111111111, 21'b000000000000010110010, 21'b000000000000001000110}, 
{21'b111111111111111111110, 21'b000000000000100100011, 21'b111111111111001101110, 21'b000000000000010100110, 21'b000000000000010001011}, 
{21'b000000000000010100111, 21'b111111111111101010010, 21'b000000000000000000001, 21'b111111111111000100111, 21'b111111111111100000001}, 
{21'b111111111111111111111, 21'b111111111111011101111, 21'b000000000000010110110, 21'b000000000000110111000, 21'b000000000000000000000}, 
{21'b111111111111101111010, 21'b111111111111101101011, 21'b000000000000000000000, 21'b000000000001001010011, 21'b111111111111011101101}, 
{21'b000000000000010101101, 21'b000000000000011101010, 21'b111111111111010100011, 21'b111111111111111100011, 21'b000000000000001111100}, 
{21'b000000000000000000000, 21'b000000000000010101011, 21'b000000000000000001001, 21'b111111111111100101011, 21'b111111111110110000010}, 
{21'b000000000000010110101, 21'b000000000000001000001, 21'b000000000000110101101, 21'b111111111111110111000, 21'b111111111111001001001}, 
{21'b000000000000001011100, 21'b111111111111111001110, 21'b111111111111010001110, 21'b111111111111111011110, 21'b000000000001000100101}, 
{21'b111111111111000011010, 21'b111111111111100000101, 21'b111111111111100011100, 21'b000000000000110011000, 21'b000000000000000100000}, 
{21'b000000000000101100010, 21'b111111111111101010000, 21'b111111111111101110101, 21'b111111111111100011000, 21'b111111111111111000010}, 
{21'b000000000000011000111, 21'b111111111111111010110, 21'b111111111111001011001, 21'b111111111111111100000, 21'b000000000000001001000}, 
{21'b000000000000100001000, 21'b000000000000000101010, 21'b111111111111100100000, 21'b000000000000000000000, 21'b111111111111001111111}, 
{21'b000000000000011101100, 21'b111111111111110100111, 21'b111111111111100100110, 21'b000000000000011010100, 21'b000000000000001100001}, 
{21'b000000000000001000101, 21'b111111111111111100000, 21'b000000000000100110000, 21'b111111111111001000110, 21'b111111111111111101010}, 
{21'b000000000000000000000, 21'b000000000000001111000, 21'b000000000000111110010, 21'b111111111110111101101, 21'b111111111110110000111}, 
{21'b111111111111110011011, 21'b000000000000001110000, 21'b000000000000010110101, 21'b111111111111010010010, 21'b000000000001000010110}, 
{21'b111111111111111111111, 21'b000000000000010101000, 21'b000000000000100100001, 21'b000000000000000100110, 21'b111111111110110110110}, 
{21'b111111111111101010010, 21'b000000000000101110101, 21'b111111111111100011011, 21'b000000000000000000101, 21'b000000000000110001101}, 
{21'b000000000000000011010, 21'b000000000000100010000, 21'b000000000000000011110, 21'b111111111110100000010, 21'b000000000001000110001}, 
{21'b111111111111000101001, 21'b111111111111100000110, 21'b000000000000011011011, 21'b000000000000011111010, 21'b000000000000011001110}, 
{21'b000000000000000000100, 21'b000000000000011110110, 21'b111111111111111011010, 21'b111111111111101100101, 21'b000000000000000100000}, 
{21'b111111111111110010101, 21'b000000000000011111100, 21'b111111111110111111100, 21'b000000000000010001110, 21'b111111111111101011101}, 
{21'b111111111111111101101, 21'b000000000000010010000, 21'b111111111111101010011, 21'b111111111111001100101, 21'b000000000001001011111}, 
{21'b000000000000111001011, 21'b000000000000001000111, 21'b000000000000101001100, 21'b111111111110110100100, 21'b111111111111010111101}, 
{21'b111111111111111000011, 21'b111111111111001110100, 21'b000000000000101110110, 21'b000000000000001001000, 21'b000000000000010000010}
};

localparam logic signed [20:0] bias [5] = '{
21'b111111111111111000000,  // -0.06223141402006149
21'b111111111111110111111,  // -0.06270556896924973
21'b111111111111110111000,  // -0.07014333456754684
21'b000000000000001010100,  // 0.0820775106549263
21'b000000000000011011100   // 0.2155742198228836
};
endpackage