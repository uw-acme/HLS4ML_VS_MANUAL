// Width: 27
// NFRAC: 13
package dense_4_27_13;

localparam logic signed [26:0] weights [32][5] = '{ 
{27'b111111111111111111110011110, 27'b000000000000000101000011001, 27'b111111111111111011001110111, 27'b000000000000000001000011011, 27'b111111111111111110010011001}, 
{27'b111111111111110111000100111, 27'b111111111111111111000111101, 27'b000000000000000111010111010, 27'b111111111111111111110011011, 27'b000000000000000000010001001}, 
{27'b000000000000000101111100011, 27'b000000000000000011011000110, 27'b111111111111111111100011010, 27'b111111111111111001100000111, 27'b111111111111111100101000000}, 
{27'b111111111111111001111111011, 27'b111111111111111010000010001, 27'b111111111111111110001101100, 27'b000000000000000100111011001, 27'b000000000000000011110000101}, 
{27'b000000000000000001111101000, 27'b000000000000000010000011110, 27'b000000000000000010100000110, 27'b111111111111111111101101010, 27'b111111111111101111110010110}, 
{27'b000000000000000101001110111, 27'b111111111111111001101100001, 27'b000000000000000010111001110, 27'b111111111111111101011010111, 27'b111111111111111101010001100}, 
{27'b111111111111111001100101000, 27'b000000000000000000100100011, 27'b111111111111111111111111111, 27'b000000000000000010110010010, 27'b000000000000000001000110101}, 
{27'b111111111111111111111110000, 27'b000000000000000100100011010, 27'b111111111111111001101110101, 27'b000000000000000010100110100, 27'b000000000000000010001011011}, 
{27'b000000000000000010100111010, 27'b111111111111111101010010100, 27'b000000000000000000000001010, 27'b111111111111111000100111011, 27'b111111111111111100000001010}, 
{27'b111111111111111111111111110, 27'b111111111111111011101111010, 27'b000000000000000010110110001, 27'b000000000000000110111000010, 27'b000000000000000000000000000}, 
{27'b111111111111111101111010111, 27'b111111111111111101101011111, 27'b000000000000000000000000000, 27'b000000000000001001010011010, 27'b111111111111111011101101111}, 
{27'b000000000000000010101101011, 27'b000000000000000011101010101, 27'b111111111111111010100011110, 27'b111111111111111111100011110, 27'b000000000000000001111100101}, 
{27'b000000000000000000000000000, 27'b000000000000000010101011101, 27'b000000000000000000001001001, 27'b111111111111111100101011001, 27'b111111111111110110000010001}, 
{27'b000000000000000010110101100, 27'b000000000000000001000001010, 27'b000000000000000110101101100, 27'b111111111111111110111000010, 27'b111111111111111001001001111}, 
{27'b000000000000000001011100111, 27'b111111111111111111001110101, 27'b111111111111111010001110111, 27'b111111111111111111011110001, 27'b000000000000001000100101001}, 
{27'b111111111111111000011010100, 27'b111111111111111100000101110, 27'b111111111111111100011100001, 27'b000000000000000110011000011, 27'b000000000000000000100000110}, 
{27'b000000000000000101100010000, 27'b111111111111111101010000001, 27'b111111111111111101110101000, 27'b111111111111111100011000111, 27'b111111111111111111000010101}, 
{27'b000000000000000011000111101, 27'b111111111111111111010110100, 27'b111111111111111001011001110, 27'b111111111111111111100000101, 27'b000000000000000001001000011}, 
{27'b000000000000000100001000101, 27'b000000000000000000101010100, 27'b111111111111111100100000110, 27'b000000000000000000000000000, 27'b111111111111111001111111001}, 
{27'b000000000000000011101100111, 27'b111111111111111110100111011, 27'b111111111111111100100110000, 27'b000000000000000011010100001, 27'b000000000000000001100001011}, 
{27'b000000000000000001000101010, 27'b111111111111111111100000111, 27'b000000000000000100110000101, 27'b111111111111111001000110101, 27'b111111111111111111101010001}, 
{27'b000000000000000000000000000, 27'b000000000000000001111000101, 27'b000000000000000111110010010, 27'b111111111111110111101101010, 27'b111111111111110110000111100}, 
{27'b111111111111111110011011011, 27'b000000000000000001110000010, 27'b000000000000000010110101011, 27'b111111111111111010010010100, 27'b000000000000001000010110111}, 
{27'b111111111111111111111111100, 27'b000000000000000010101000110, 27'b000000000000000100100001011, 27'b000000000000000000100110111, 27'b111111111111110110110110001}, 
{27'b111111111111111101010010101, 27'b000000000000000101110101000, 27'b111111111111111100011011000, 27'b000000000000000000000101110, 27'b000000000000000110001101011}, 
{27'b000000000000000000011010111, 27'b000000000000000100010000000, 27'b000000000000000000011110010, 27'b111111111111110100000010000, 27'b000000000000001000110001011}, 
{27'b111111111111111000101001010, 27'b111111111111111100000110100, 27'b000000000000000011011011010, 27'b000000000000000011111010011, 27'b000000000000000011001110100}, 
{27'b000000000000000000000100001, 27'b000000000000000011110110110, 27'b111111111111111111011010100, 27'b111111111111111101100101111, 27'b000000000000000000100000011}, 
{27'b111111111111111110010101010, 27'b000000000000000011111100000, 27'b111111111111110111111100000, 27'b000000000000000010001110000, 27'b111111111111111101011101110}, 
{27'b111111111111111111101101001, 27'b000000000000000010010000100, 27'b111111111111111101010011001, 27'b111111111111111001100101111, 27'b000000000000001001011111110}, 
{27'b000000000000000111001011101, 27'b000000000000000001000111100, 27'b000000000000000101001100010, 27'b111111111111110110100100000, 27'b111111111111111010111101010}, 
{27'b111111111111111111000011011, 27'b111111111111111001110100100, 27'b000000000000000101110110100, 27'b000000000000000001001000100, 27'b000000000000000010000010100}
};

localparam logic signed [26:0] bias [5] = '{
27'b111111111111111111000000010,  // -0.06223141402006149
27'b111111111111111110111111110,  // -0.06270556896924973
27'b111111111111111110111000001,  // -0.07014333456754684
27'b000000000000000001010100000,  // 0.0820775106549263
27'b000000000000000011011100101   // 0.2155742198228836
};
endpackage