// Width: 19
// NFRAC: 9
package dense_1_19_9;

localparam logic signed [18:0] weights [16][64] = '{ 
{19'b0000000000010000010, 19'b1111111111010110010, 19'b1111111111110100011, 19'b1111111111110001100, 19'b1111111111100110000, 19'b0000000000000111000, 19'b1111111110111101101, 19'b0000000000000000000, 19'b0000000000000011101, 19'b0000000000010000110, 19'b0000000000000000001, 19'b1111111111100110000, 19'b1111111111111111111, 19'b0000000000001101011, 19'b0000000000000010001, 19'b1111111111101111010, 19'b0000000000001110111, 19'b0000000000000011110, 19'b0000000000000000000, 19'b1111111111111111111, 19'b0000000000011000000, 19'b1111111111101010110, 19'b1111111111111110100, 19'b0000000000011110010, 19'b1111111111101011011, 19'b1111111111010100010, 19'b1111111111101110010, 19'b1111111111110011100, 19'b1111111111111001010, 19'b1111111111111111111, 19'b0000000000000010011, 19'b0000000000001111101, 19'b0000000000001100100, 19'b1111111111111111001, 19'b0000000000000000000, 19'b0000000000010011111, 19'b1111111111111110110, 19'b1111111111101111111, 19'b0000000000000001101, 19'b0000000000001100010, 19'b1111111111111111001, 19'b0000000000010001100, 19'b1111111111101110111, 19'b0000000000111011011, 19'b1111111111111111111, 19'b0000000000011100111, 19'b0000000000000000000, 19'b0000000000001011110, 19'b0000000000001100100, 19'b1111111111111110011, 19'b0000000000000000000, 19'b0000000000001010010, 19'b0000000000001101110, 19'b0000000000000100111, 19'b1111111111111000100, 19'b1111111111101100001, 19'b0000000000100010010, 19'b1111111111100000000, 19'b0000000000011101111, 19'b1111111111101001010, 19'b0000000000110010110, 19'b1111111111111111100, 19'b0000000000000000101, 19'b0000000000000101001}, 
{19'b0000000000000000001, 19'b1111111111101011011, 19'b1111111111110111100, 19'b1111111111101110000, 19'b1111111111101011101, 19'b0000000000000110110, 19'b1111111111001111101, 19'b1111111111111111110, 19'b1111111111110001011, 19'b0000000000001011000, 19'b0000000000000000011, 19'b1111111111111010011, 19'b0000000000001100100, 19'b0000000000000000000, 19'b1111111111111111111, 19'b0000000000001101010, 19'b1111111111111111100, 19'b0000000000000000000, 19'b1111111111110100010, 19'b1111111111101111111, 19'b0000000000011100010, 19'b1111111111111010110, 19'b0000000000000011000, 19'b0000000000101100101, 19'b0000000000010000011, 19'b1111111111110001010, 19'b1111111111110001001, 19'b1111111111111111111, 19'b1111111111111001100, 19'b1111111111100110000, 19'b1111111111111100001, 19'b0000000000011101000, 19'b0000000000010001110, 19'b0000000000100011001, 19'b0000000000101000010, 19'b0000000000000011001, 19'b1111111111111000011, 19'b1111111111100100001, 19'b0000000000000011101, 19'b0000000000001100000, 19'b0000000000000001011, 19'b0000000000001101001, 19'b1111111111110010011, 19'b0000000000010000001, 19'b0000000000001011000, 19'b0000000000000011001, 19'b1111111111101010001, 19'b0000000000000101000, 19'b0000000000010000101, 19'b0000000000000001111, 19'b0000000000000001100, 19'b0000000001001010000, 19'b1111111111111011001, 19'b1111111111111001101, 19'b1111111111111100100, 19'b1111111111111111100, 19'b0000000000010000011, 19'b1111111111101000010, 19'b0000000000111111000, 19'b0000000000000000010, 19'b0000000000100001010, 19'b0000000000001111010, 19'b0000000000110100101, 19'b0000000000001001000}, 
{19'b1111111111111111100, 19'b0000000000000000000, 19'b1111111111111010101, 19'b1111111111110100101, 19'b1111111111110100001, 19'b0000000000000010101, 19'b0000000001011110110, 19'b1111111111111111111, 19'b1111111110101110111, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111111110110, 19'b1111111111110001011, 19'b0000000000000000000, 19'b1111111111111111011, 19'b0000000000001010110, 19'b0000000000111001111, 19'b1111111111111111111, 19'b0000000000000100100, 19'b0000000000000000000, 19'b0000000000011010011, 19'b1111111111010001110, 19'b0000000000100100111, 19'b1111111111010010010, 19'b0000000000111100101, 19'b1111111111101001110, 19'b1111111111110000010, 19'b1111111111010010000, 19'b0000000001010001100, 19'b0000000000010001101, 19'b0000000000000000101, 19'b0000000000100001001, 19'b0000000001000001010, 19'b1111111110110011100, 19'b1111111111111001111, 19'b0000000000000010000, 19'b1111111111110001001, 19'b0000000000111001011, 19'b1111111111111101011, 19'b0000000000010100000, 19'b0000000000010101010, 19'b0000000000010111101, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111111110111, 19'b0000000000001010000, 19'b1111111111101110000, 19'b1111111111110101000, 19'b1111111111111110111, 19'b0000000000011001001, 19'b1111111111110100101, 19'b0000000000001001100, 19'b1111111111111111111, 19'b0000000000001000100, 19'b1111111111110100110, 19'b1111111111111111111, 19'b1111111111101100010, 19'b1111111111010101001, 19'b1111111111111111110, 19'b0000000000000000000, 19'b0000000001100010101, 19'b0000000000000000110, 19'b1111111111111111110, 19'b1111111111101100001}, 
{19'b1111111111100010101, 19'b1111111111101000011, 19'b1111111111010011101, 19'b0000000000010011101, 19'b1111111111101011110, 19'b1111111110101001110, 19'b1111111111111000101, 19'b1111111111101100010, 19'b0000000000001110010, 19'b1111111111111111111, 19'b0000000001010000111, 19'b1111111111111001001, 19'b1111111111001101111, 19'b0000000000100101000, 19'b0000000000000001100, 19'b1111111111111111111, 19'b1111111111100011100, 19'b1111111111111111111, 19'b0000000000000000000, 19'b1111111111110001100, 19'b1111111110110110010, 19'b1111111111111000110, 19'b1111111111010011010, 19'b0000000000001100101, 19'b1111111111100111001, 19'b1111111111000101000, 19'b0000000000010100000, 19'b0000000000101111001, 19'b0000000001010010111, 19'b1111111111100010100, 19'b1111111111011010101, 19'b0000000000000100101, 19'b0000000000100000000, 19'b1111111111001010001, 19'b1111111111101011111, 19'b0000000000000000000, 19'b1111111111010001100, 19'b0000000000001111100, 19'b1111111111100011110, 19'b0000000000000111101, 19'b0000000000011101010, 19'b0000000000001010000, 19'b0000000000000000000, 19'b0000000000000001010, 19'b0000000000100011010, 19'b1111111111110011001, 19'b1111111111111111111, 19'b1111111111101001111, 19'b1111111111111111111, 19'b1111111111111001110, 19'b1111111111011000100, 19'b0000000000000101100, 19'b1111111111111111111, 19'b0000000000001101111, 19'b0000000000010100001, 19'b0000000000101001011, 19'b1111111111000010000, 19'b1111111111000100100, 19'b1111111111010010110, 19'b0000000000110111011, 19'b0000000001101111111, 19'b1111111111000110011, 19'b1111111111111100100, 19'b0000000000011011110}, 
{19'b0000000000010101111, 19'b1111111111011000011, 19'b1111111111101111011, 19'b1111111111111111111, 19'b1111111111110110001, 19'b0000000000010101110, 19'b0000000000001100001, 19'b1111111111111111111, 19'b1111111111011001110, 19'b1111111111110000100, 19'b1111111111101000011, 19'b0000000000000011011, 19'b0000000000000000000, 19'b0000000000000000000, 19'b1111111111111101011, 19'b0000000000010110111, 19'b0000000000001000100, 19'b1111111111100110110, 19'b0000000000000001111, 19'b0000000000000000110, 19'b0000000000001101011, 19'b1111111111111000011, 19'b0000000000000100110, 19'b1111111111111110110, 19'b0000000001000100001, 19'b1111111111110100000, 19'b1111111111101110000, 19'b1111111111100110001, 19'b0000000000000000000, 19'b0000000000001010100, 19'b0000000000000111011, 19'b0000000000010001100, 19'b1111111111111111001, 19'b0000000000000100101, 19'b0000000000001000010, 19'b1111111111111111111, 19'b0000000000000000011, 19'b0000000000111000011, 19'b1111111111101101100, 19'b1111111111111011000, 19'b0000000000011011101, 19'b0000000000001111111, 19'b1111111111100000101, 19'b0000000000000000011, 19'b1111111110111011101, 19'b1111111111111111111, 19'b1111111111111000001, 19'b0000000000000000110, 19'b1111111111111111111, 19'b1111111111111110011, 19'b1111111111111111111, 19'b0000000000001100000, 19'b1111111111111111101, 19'b0000000000010100010, 19'b1111111111110011110, 19'b1111111111010000111, 19'b1111111111100010001, 19'b1111111111011111011, 19'b1111111111011000101, 19'b0000000000101111110, 19'b0000000001010111111, 19'b0000000000110010101, 19'b0000000000000111110, 19'b1111111111111111111}, 
{19'b1111111111100011011, 19'b1111111111010111101, 19'b0000000000000000000, 19'b0000000000010011101, 19'b0000000000010010010, 19'b1111111111110010011, 19'b0000000000100101010, 19'b1111111111111111111, 19'b0000000000001111100, 19'b1111111111111111111, 19'b1111111111111111011, 19'b1111111111111011010, 19'b1111111111110100101, 19'b0000000000100101000, 19'b1111111111111010010, 19'b0000000000000000000, 19'b1111111111011000000, 19'b1111111111101001010, 19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111111111100111, 19'b1111111111101011111, 19'b1111111111101011100, 19'b0000000000011101110, 19'b1111111111101011101, 19'b1111111111111111111, 19'b0000000000010000011, 19'b1111111111111011010, 19'b1111111111000100010, 19'b1111111111111111111, 19'b1111111111111011101, 19'b1111111111111111010, 19'b1111111111111111010, 19'b0000000000000010100, 19'b0000000000001000011, 19'b0000000000010110001, 19'b0000000000000000110, 19'b1111111111111001101, 19'b1111111111101111001, 19'b1111111111111111111, 19'b1111111111110101001, 19'b1111111111011110011, 19'b0000000000011001100, 19'b0000000000000000101, 19'b0000000000100110100, 19'b0000000000000000000, 19'b1111111111111111111, 19'b0000000000000110000, 19'b1111111111100101001, 19'b0000000000001110111, 19'b0000000000000000000, 19'b1111111111111001100, 19'b1111111111101000110, 19'b0000000000011000101, 19'b1111111111111111111, 19'b0000000000010110001, 19'b0000000000001101110, 19'b0000000000001101000, 19'b1111111111111110110, 19'b1111111111111111011, 19'b1111111111001100010, 19'b1111111111110111111, 19'b1111111111111100010, 19'b1111111111111111111}, 
{19'b1111111111101101111, 19'b1111111111101010100, 19'b1111111111100100011, 19'b1111111111111011100, 19'b1111111111110111011, 19'b0000000000000110101, 19'b1111111111010011010, 19'b1111111111110110011, 19'b1111111111110001101, 19'b1111111111111111111, 19'b1111111111101101100, 19'b0000000000010110010, 19'b0000000000000010010, 19'b0000000000001000110, 19'b0000000000010011111, 19'b0000000000000000000, 19'b0000000000110011000, 19'b0000000000000101101, 19'b0000000000001111100, 19'b0000000000010001001, 19'b1111111111110101111, 19'b0000000000010111010, 19'b1111111111110000011, 19'b1111111111011111111, 19'b0000000000001011000, 19'b0000000000100001000, 19'b1111111111111111101, 19'b0000000000000011011, 19'b1111111111000011001, 19'b0000000000010010010, 19'b0000000000010001000, 19'b1111111111101000000, 19'b0000000000011110001, 19'b0000000000101010100, 19'b0000000000000000000, 19'b0000000000010101111, 19'b1111111111111111111, 19'b0000000000010010001, 19'b0000000000001100101, 19'b0000000000000000000, 19'b1111111111111000011, 19'b1111111111101000101, 19'b0000000000001001001, 19'b0000000000011110111, 19'b0000000000100001001, 19'b1111111111110101001, 19'b1111111111111010101, 19'b1111111111110011110, 19'b1111111111110111010, 19'b0000000000000111100, 19'b0000000000000000001, 19'b0000000000000010001, 19'b0000000000000000000, 19'b0000000000001011100, 19'b1111111111110100110, 19'b0000000000110001010, 19'b0000000000010110110, 19'b1111111111111110011, 19'b0000000000011000111, 19'b0000000000001101111, 19'b1111111110010111111, 19'b1111111111011011000, 19'b1111111111110100111, 19'b1111111111111111010}, 
{19'b0000000000000000010, 19'b0000000000001111010, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111101011011, 19'b1111111111111110000, 19'b1111111111101111100, 19'b0000000000000000000, 19'b0000000000000001110, 19'b0000000000011000111, 19'b0000000000000000111, 19'b1111111111100111110, 19'b1111111111111011111, 19'b0000000000000000000, 19'b1111111111111100101, 19'b1111111111100011001, 19'b1111111111001001101, 19'b1111111111111111111, 19'b1111111111011001010, 19'b1111111111100011011, 19'b1111111111100111000, 19'b0000000000010110001, 19'b0000000000000011000, 19'b1111111111110110111, 19'b1111111111100100000, 19'b0000000000001001111, 19'b0000000000000000000, 19'b0000000000011111111, 19'b0000000000110011100, 19'b1111111111111101011, 19'b0000000000000000000, 19'b0000000000001110110, 19'b1111111111010100010, 19'b1111111111101000010, 19'b0000000000000011100, 19'b0000000000000101111, 19'b1111111111101110000, 19'b0000000000001111010, 19'b0000000000001000011, 19'b1111111111110110001, 19'b1111111111100101001, 19'b1111111111111101101, 19'b0000000000000010000, 19'b1111111111110101010, 19'b0000000000000011100, 19'b0000000000001110101, 19'b1111111111111000010, 19'b0000000000000001100, 19'b0000000000000000000, 19'b1111111111110010000, 19'b1111111111100111001, 19'b0000000000011010100, 19'b0000000000001000000, 19'b1111111111110100100, 19'b0000000000001000011, 19'b1111111111111100000, 19'b1111111111100001101, 19'b1111111111110111011, 19'b1111111111111100101, 19'b1111111111111011100, 19'b0000000000110101001, 19'b0000000000001100001, 19'b1111111111111100111, 19'b1111111111111111111}, 
{19'b0000000000000000111, 19'b0000000000100101100, 19'b1111111111011010110, 19'b1111111111110001001, 19'b0000000000010100101, 19'b1111111111110010110, 19'b0000000001001101100, 19'b1111111111101101100, 19'b1111111111111111111, 19'b0000000000010010110, 19'b0000000000010000010, 19'b1111111111111111110, 19'b1111111111111100111, 19'b1111111111100001001, 19'b0000000000010010000, 19'b0000000000001010001, 19'b1111111111110011100, 19'b1111111111111111111, 19'b0000000000000000000, 19'b0000000000000000000, 19'b0000000000010000111, 19'b1111111111100010100, 19'b0000000000011001000, 19'b0000000000100111001, 19'b1111111111111010011, 19'b1111111111111111111, 19'b1111111111111110111, 19'b1111111111111111111, 19'b0000000000101111000, 19'b0000000000000000010, 19'b1111111111101110100, 19'b0000000000000000000, 19'b0000000000011000100, 19'b1111111111001100000, 19'b1111111111011101011, 19'b0000000000001100101, 19'b0000000000001000110, 19'b1111111111011011011, 19'b1111111111110011111, 19'b1111111111110010010, 19'b0000000000011001101, 19'b0000000000011001000, 19'b0000000000000000000, 19'b1111111111101110101, 19'b0000000000000000000, 19'b0000000000011001010, 19'b1111111111111100001, 19'b1111111111111111111, 19'b0000000000000000101, 19'b0000000000001111101, 19'b1111111111111100010, 19'b1111111111110011100, 19'b0000000000010110000, 19'b1111111111110010001, 19'b0000000000010001111, 19'b0000000000100101011, 19'b0000000000000010100, 19'b0000000000010000110, 19'b1111111111100110011, 19'b1111111111101000100, 19'b0000000000110101001, 19'b1111111111110111110, 19'b0000000000000010111, 19'b1111111111111010000}, 
{19'b0000000000000001000, 19'b1111111111100011000, 19'b0000000000010111100, 19'b1111111111101101110, 19'b1111111111111111110, 19'b0000000000001101100, 19'b1111111111011010110, 19'b0000000000001100010, 19'b0000000000011111011, 19'b0000000000001001110, 19'b0000000000010111001, 19'b0000000000010100101, 19'b1111111111101100011, 19'b1111111111111011001, 19'b1111111111111100101, 19'b0000000000000000000, 19'b1111111111000010100, 19'b0000000000010100101, 19'b1111111111111101101, 19'b0000000000000001111, 19'b1111111111101001011, 19'b0000000000000100011, 19'b0000000000001001110, 19'b1111111111111111111, 19'b1111111111100010100, 19'b1111111111111100111, 19'b1111111111111010110, 19'b0000000001001111110, 19'b1111111111010101100, 19'b0000000000000100010, 19'b0000000000000110001, 19'b1111111111111100010, 19'b1111111111110001110, 19'b0000000000000111011, 19'b1111111111111010111, 19'b1111111111110111011, 19'b1111111111110100100, 19'b1111111111110010100, 19'b1111111111111110100, 19'b1111111111101100111, 19'b0000000000010100100, 19'b0000000000000111111, 19'b0000000000011111110, 19'b0000000000000101100, 19'b0000000000000010010, 19'b1111111111101101011, 19'b0000000000000000000, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000001100011, 19'b0000000000001011010, 19'b0000000000010010110, 19'b1111111111111111100, 19'b1111111111101101001, 19'b0000000000000000100, 19'b0000000000000000000, 19'b0000000000010100101, 19'b1111111111110011001, 19'b1111111111011100110, 19'b0000000000100011111, 19'b1111111111101101001, 19'b0000000001001010011, 19'b1111111111111110101, 19'b1111111111101001010}, 
{19'b1111111111011011000, 19'b1111111111111111111, 19'b1111111111100101110, 19'b0000000000001110101, 19'b0000000000010000110, 19'b1111111111111001011, 19'b0000000000100001000, 19'b1111111111110101000, 19'b1111111111100001010, 19'b1111111111101000100, 19'b1111111111101111111, 19'b1111111111100001100, 19'b1111111111110001010, 19'b0000000000001100100, 19'b0000000000000000000, 19'b0000000000000000000, 19'b0000000000110101111, 19'b1111111111111101001, 19'b1111111111111111111, 19'b0000000000011010010, 19'b0000000000010010101, 19'b1111111111011010111, 19'b1111111111100111100, 19'b0000000000001100000, 19'b1111111111100100011, 19'b1111111111111110101, 19'b1111111111101111011, 19'b1111111111101010100, 19'b1111111111100100000, 19'b0000000000010011010, 19'b0000000000001110100, 19'b1111111111110110000, 19'b1111111111111011010, 19'b1111111111000001101, 19'b1111111111110100101, 19'b0000000000000011001, 19'b1111111111110111101, 19'b1111111111101101000, 19'b1111111111111111110, 19'b0000000000000111100, 19'b1111111111111000011, 19'b1111111111111111110, 19'b1111111111111101110, 19'b1111111111010101011, 19'b0000000000000000000, 19'b0000000000000000000, 19'b0000000000010101110, 19'b1111111111111000000, 19'b0000000000011011000, 19'b1111111111110011110, 19'b0000000000010010011, 19'b1111111111111111111, 19'b0000000000001110011, 19'b1111111111100110111, 19'b1111111111111111111, 19'b0000000000100000110, 19'b0000000000010100000, 19'b0000000000010010101, 19'b0000000000000001100, 19'b1111111111100110011, 19'b1111111111101100110, 19'b1111111111010100000, 19'b1111111111111111111, 19'b0000000000000110110}, 
{19'b0000000000010011101, 19'b0000000000000000001, 19'b0000000000001000011, 19'b1111111111111111111, 19'b0000000000001001110, 19'b1111111111110111011, 19'b0000000000001111000, 19'b0000000000000010101, 19'b0000000000001000101, 19'b0000000000010101110, 19'b1111111111101111001, 19'b1111111111111110101, 19'b1111111111111111011, 19'b1111111111111111011, 19'b1111111111010101110, 19'b1111111111101100111, 19'b0000000000101000010, 19'b1111111111111110001, 19'b1111111111111100101, 19'b0000000000000000000, 19'b1111111111100111101, 19'b0000000000000000100, 19'b0000000000010000000, 19'b0000000000000010011, 19'b0000000000000010010, 19'b0000000000010101101, 19'b0000000000000000000, 19'b0000000000000010011, 19'b0000000000000000000, 19'b1111111111111100111, 19'b1111111111110011001, 19'b1111111111010101011, 19'b0000000000010000111, 19'b0000000000010101111, 19'b1111111111111110001, 19'b1111111111110000111, 19'b0000000000000000000, 19'b1111111111010110000, 19'b1111111111111101000, 19'b1111111111111111110, 19'b0000000000001100100, 19'b1111111111110111101, 19'b1111111111111111111, 19'b0000000000110110001, 19'b0000000000011100101, 19'b1111111111111111100, 19'b1111111111111111111, 19'b1111111111111111111, 19'b1111111111110000100, 19'b0000000000001001011, 19'b0000000000001001001, 19'b0000000000001011001, 19'b0000000000001010000, 19'b0000000000011000110, 19'b0000000000010110011, 19'b0000000000101010001, 19'b1111111111110111000, 19'b0000000000011001001, 19'b0000000000001001110, 19'b1111111111101011001, 19'b0000000000000111000, 19'b1111111111100111001, 19'b1111111111100011110, 19'b1111111111100000000}, 
{19'b0000000000000000000, 19'b0000000000001110100, 19'b1111111111110011100, 19'b0000000000000000000, 19'b1111111111111100110, 19'b1111111111111101110, 19'b1111111111010101101, 19'b1111111111111111111, 19'b0000000000010000001, 19'b0000000000001111111, 19'b0000000000001111001, 19'b1111111111100110100, 19'b1111111111111010010, 19'b0000000000010010001, 19'b1111111111111111111, 19'b0000000000000000010, 19'b1111111111001010001, 19'b1111111111111111111, 19'b0000000000010111110, 19'b0000000000000100100, 19'b0000000000001111001, 19'b1111111111111000100, 19'b0000000000001111111, 19'b0000000000011001111, 19'b1111111111101001010, 19'b1111111111101110000, 19'b1111111111111111101, 19'b1111111111111010110, 19'b0000000000000100010, 19'b0000000000000000000, 19'b1111111111111111111, 19'b0000000000010100000, 19'b1111111111010000000, 19'b0000000000010111001, 19'b0000000000100000000, 19'b0000000000000111011, 19'b0000000000000111001, 19'b1111111111111001000, 19'b0000000000000111010, 19'b1111111111111001001, 19'b1111111111101111111, 19'b1111111111111100110, 19'b0000000000001010100, 19'b0000000000101100110, 19'b1111111111001001110, 19'b1111111111100011011, 19'b0000000000001100010, 19'b1111111111111001101, 19'b0000000000011100110, 19'b1111111111110000111, 19'b1111111111101010110, 19'b1111111111101110000, 19'b1111111111111111111, 19'b0000000000000111101, 19'b1111111111110101111, 19'b1111111111001010011, 19'b1111111111110110110, 19'b1111111111111111010, 19'b0000000000000010110, 19'b1111111111011000111, 19'b0000000001000111101, 19'b1111111111011101001, 19'b0000000000100010101, 19'b0000000000001001110}, 
{19'b0000000000000101000, 19'b1111111111110011101, 19'b0000000000101000001, 19'b1111111111101100101, 19'b1111111111100010010, 19'b0000000000000101110, 19'b0000000000010011110, 19'b0000000000010011001, 19'b1111111111110100101, 19'b1111111111110101101, 19'b0000000000000011010, 19'b0000000000001110101, 19'b0000000000001111000, 19'b0000000000000011001, 19'b1111111111110010111, 19'b0000000000001000001, 19'b0000000000011110001, 19'b1111111111111111010, 19'b1111111111101110000, 19'b0000000000000000000, 19'b0000000000000100110, 19'b0000000000000001010, 19'b1111111111101101001, 19'b0000000000000111001, 19'b0000000000110010010, 19'b0000000000000000101, 19'b0000000000001011100, 19'b1111111111001101001, 19'b1111111111111011010, 19'b0000000000000000100, 19'b1111111111110011011, 19'b1111111111101100000, 19'b0000000000011101010, 19'b1111111111111110010, 19'b1111111111111101100, 19'b1111111111101100011, 19'b0000000000001000110, 19'b0000000000010010101, 19'b1111111111111111011, 19'b1111111111111101001, 19'b1111111111110100000, 19'b0000000000001110100, 19'b0000000000000000000, 19'b1111111111010100000, 19'b0000000000010011111, 19'b0000000000011001100, 19'b1111111111111111111, 19'b0000000000000001101, 19'b1111111111100100001, 19'b1111111111111011001, 19'b1111111111111111111, 19'b1111111111101011101, 19'b0000000000000000000, 19'b1111111111110100111, 19'b0000000000000011101, 19'b1111111111001011101, 19'b1111111111111111111, 19'b1111111111111111111, 19'b0000000000010001100, 19'b0000000000100100000, 19'b1111111111010011100, 19'b0000000000100001010, 19'b0000000000000010010, 19'b1111111111111011001}, 
{19'b0000000000010010011, 19'b0000000001001111011, 19'b0000000000011111101, 19'b0000000000010010010, 19'b1111111111100001011, 19'b1111111111101011101, 19'b1111111101011001101, 19'b1111111111100010110, 19'b0000000000011001110, 19'b1111111111111111111, 19'b0000000000010010110, 19'b0000000000110111001, 19'b0000000000000100011, 19'b0000000000000000010, 19'b1111111111111110111, 19'b0000000000000000000, 19'b1111111111110011111, 19'b1111111111110011000, 19'b0000000000001110101, 19'b1111111111011111110, 19'b1111111111010101011, 19'b1111111111111001011, 19'b1111111111011010101, 19'b0000000000000001111, 19'b1111111101101110010, 19'b0000000000110100001, 19'b0000000000111111010, 19'b0000000000100110101, 19'b1111111110010000011, 19'b1111111111101011111, 19'b1111111111010011111, 19'b1111111111001010000, 19'b1111111101011110011, 19'b0000000000101011010, 19'b1111111111111101001, 19'b0000000000010100011, 19'b0000000000000001100, 19'b1111111110100100010, 19'b0000000000000000000, 19'b0000000000000000000, 19'b0000000000000010000, 19'b0000000001000001001, 19'b1111111111110010111, 19'b1111111111010110101, 19'b0000000000111001011, 19'b1111111111100011100, 19'b1111111111101011001, 19'b1111111111100110111, 19'b0000000000011110100, 19'b0000000000100010000, 19'b1111111111111011101, 19'b1111111111101001101, 19'b1111111111111111110, 19'b1111111111111000110, 19'b0000000000000000000, 19'b1111111111100111110, 19'b0000000000100110110, 19'b0000000001000101011, 19'b0000000000101101100, 19'b1111111111000101110, 19'b1111111100010011000, 19'b0000000000111000101, 19'b0000000000000101111, 19'b0000000000010100010}, 
{19'b1111111111110000100, 19'b0000000000010101100, 19'b0000000000010100010, 19'b1111111111111111111, 19'b1111111111101000001, 19'b1111111111111010010, 19'b1111111111100111011, 19'b1111111111111100011, 19'b0000000000001001100, 19'b1111111111111011001, 19'b1111111111111110000, 19'b1111111111111101011, 19'b1111111111111111111, 19'b1111111111110100010, 19'b1111111111111110010, 19'b1111111111111001100, 19'b0000000000010100000, 19'b1111111111111111111, 19'b1111111111010110111, 19'b0000000000011101110, 19'b0000000000100110000, 19'b0000000000011010100, 19'b1111111111101011101, 19'b1111111111110111001, 19'b1111111111101001110, 19'b1111111111101101011, 19'b0000000000001110100, 19'b0000000000001110111, 19'b0000000000001110011, 19'b0000000000010111000, 19'b0000000000000010001, 19'b0000000000011000101, 19'b1111111111111101010, 19'b0000000000000000010, 19'b0000000000010011011, 19'b0000000000001000011, 19'b1111111111111011110, 19'b1111111111111111011, 19'b0000000000000000000, 19'b1111111111101101010, 19'b1111111111110001101, 19'b1111111111111000111, 19'b1111111111101001000, 19'b0000000000011100110, 19'b0000000000000000000, 19'b1111111111111111101, 19'b1111111111111010101, 19'b1111111111110110100, 19'b1111111111001100011, 19'b1111111111111101100, 19'b1111111111110001101, 19'b1111111111110110111, 19'b1111111111111001100, 19'b0000000000010000111, 19'b0000000000101011101, 19'b0000000000001011111, 19'b1111111111111111001, 19'b1111111111101010000, 19'b1111111111111110000, 19'b0000000000000000000, 19'b0000000000010100110, 19'b1111111111111110101, 19'b0000000000000010111, 19'b0000000000000000000}
};

localparam logic signed [18:0] bias [64] = '{
19'b1111111111111101100,  // -0.037350185215473175
19'b0000000000010001100,  // 0.27355897426605225
19'b1111111111111000000,  // -0.12378914654254913
19'b1111111111111011110,  // -0.064457006752491
19'b0000000000000011011,  // 0.05452875792980194
19'b0000000000000111011,  // 0.11671770364046097
19'b0000000000001000101,  // 0.13640816509723663
19'b0000000000000100110,  // 0.07482525706291199
19'b0000000000000010111,  // 0.04674031585454941
19'b1111111111110011000,  // -0.20146161317825317
19'b1111111111111001101,  // -0.09910125285387039
19'b0000000000001001101,  // 0.15104414522647858
19'b1111111111111001011,  // -0.10221704095602036
19'b1111111111110110101,  // -0.1461549550294876
19'b1111111111111010011,  // -0.08641516417264938
19'b0000000000001010101,  // 0.16613510251045227
19'b1111111111111010101,  // -0.0836295336484909
19'b1111111111111100010,  // -0.05756539851427078
19'b1111111111111101111,  // -0.03229188174009323
19'b1111111111111110001,  // -0.028388574719429016
19'b0000000000001000000,  // 0.1260243058204651
19'b1111111111111101101,  // -0.037064336240291595
19'b0000000000001100011,  // 0.19336333870887756
19'b0000000000000001010,  // 0.02124214917421341
19'b0000000000011111111,  // 0.4985624849796295
19'b0000000000000001000,  // 0.0158411655575037
19'b1111111111111010101,  // -0.08296407759189606
19'b0000000000000111000,  // 0.11056788265705109
19'b0000000000000000110,  // 0.01173810102045536
19'b1111111111111001000,  // -0.10843746364116669
19'b0000000000010001100,  // 0.27439257502555847
19'b0000000000000101111,  // 0.09199801832437515
19'b0000000000010001100,  // 0.27419957518577576
19'b0000000000010001010,  // 0.27063727378845215
19'b1111111111110000000,  // -0.24828937649726868
19'b0000000000000101000,  // 0.07818280160427094
19'b1111111111111111101,  // -0.005749030504375696
19'b0000000000000110111,  // 0.10850494354963303
19'b0000000000001000101,  // 0.13591453433036804
19'b1111111111111000010,  // -0.12088628858327866
19'b1111111111111100010,  // -0.05666546896100044
19'b0000000000000101111,  // 0.09311636537313461
19'b0000000000000011100,  // 0.05477767437696457
19'b0000000000000001111,  // 0.029585206881165504
19'b1111111111101100000,  // -0.31209176778793335
19'b1111111111111010100,  // -0.08465463668107986
19'b1111111111110101010,  // -0.16775836050510406
19'b0000000000001001011,  // 0.14762157201766968
19'b1111111111110000111,  // -0.23618532717227936
19'b0000000000000100001,  // 0.06535740196704865
19'b1111111111110111110,  // -0.12853026390075684
19'b1111111111110111001,  // -0.13802281022071838
19'b1111111111110110010,  // -0.15156887471675873
19'b0000000000000101000,  // 0.07979883998632431
19'b0000000000001011100,  // 0.18141601979732513
19'b1111111111111100100,  // -0.054039113223552704
19'b1111111111111111010,  // -0.010052933357656002
19'b0000000000000100001,  // 0.06611225008964539
19'b0000000000000011001,  // 0.05053366720676422
19'b0000000000000001101,  // 0.026860840618610382
19'b0000000000000010000,  // 0.03283466026186943
19'b0000000000001001111,  // 0.15558314323425293
19'b1111111111101101101,  // -0.2863388657569885
19'b1111111111111010011   // -0.08769102394580841
};
endpackage