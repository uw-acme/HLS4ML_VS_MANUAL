// Width: 28
// NFRAC: 14
package dense_4_28_14;

localparam logic signed [27:0] weights [32][5] = '{ 
{28'b1111111111111111111100111101, 28'b0000000000000001010000110011, 28'b1111111111111110110011101110, 28'b0000000000000000010000110110, 28'b1111111111111111100100110010}, 
{28'b1111111111111101110001001111, 28'b1111111111111111110001111011, 28'b0000000000000001110101110100, 28'b1111111111111111111100110110, 28'b0000000000000000000100010010}, 
{28'b0000000000000001011111000111, 28'b0000000000000000110110001101, 28'b1111111111111111111000110101, 28'b1111111111111110011000001110, 28'b1111111111111111001010000001}, 
{28'b1111111111111110011111110110, 28'b1111111111111110100000100010, 28'b1111111111111111100011011000, 28'b0000000000000001001110110011, 28'b0000000000000000111100001010}, 
{28'b0000000000000000011111010001, 28'b0000000000000000100000111100, 28'b0000000000000000101000001101, 28'b1111111111111111111011010100, 28'b1111111111111011111100101100}, 
{28'b0000000000000001010011101110, 28'b1111111111111110011011000010, 28'b0000000000000000101110011100, 28'b1111111111111111010110101110, 28'b1111111111111111010100011001}, 
{28'b1111111111111110011001010001, 28'b0000000000000000001001000111, 28'b1111111111111111111111111111, 28'b0000000000000000101100100101, 28'b0000000000000000010001101010}, 
{28'b1111111111111111111111100000, 28'b0000000000000001001000110101, 28'b1111111111111110011011101011, 28'b0000000000000000101001101001, 28'b0000000000000000100010110110}, 
{28'b0000000000000000101001110100, 28'b1111111111111111010100101000, 28'b0000000000000000000000010101, 28'b1111111111111110001001110111, 28'b1111111111111111000000010101}, 
{28'b1111111111111111111111111100, 28'b1111111111111110111011110101, 28'b0000000000000000101101100010, 28'b0000000000000001101110000100, 28'b0000000000000000000000000000}, 
{28'b1111111111111111011110101110, 28'b1111111111111111011010111111, 28'b0000000000000000000000000000, 28'b0000000000000010010100110101, 28'b1111111111111110111011011110}, 
{28'b0000000000000000101011010111, 28'b0000000000000000111010101010, 28'b1111111111111110101000111100, 28'b1111111111111111111000111101, 28'b0000000000000000011111001010}, 
{28'b0000000000000000000000000001, 28'b0000000000000000101010111010, 28'b0000000000000000000010010010, 28'b1111111111111111001010110011, 28'b1111111111111101100000100011}, 
{28'b0000000000000000101101011000, 28'b0000000000000000010000010101, 28'b0000000000000001101011011001, 28'b1111111111111111101110000100, 28'b1111111111111110010010011110}, 
{28'b0000000000000000010111001111, 28'b1111111111111111110011101011, 28'b1111111111111110100011101110, 28'b1111111111111111110111100011, 28'b0000000000000010001001010011}, 
{28'b1111111111111110000110101000, 28'b1111111111111111000001011101, 28'b1111111111111111000111000011, 28'b0000000000000001100110000111, 28'b0000000000000000001000001101}, 
{28'b0000000000000001011000100001, 28'b1111111111111111010100000010, 28'b1111111111111111011101010000, 28'b1111111111111111000110001111, 28'b1111111111111111110000101010}, 
{28'b0000000000000000110001111011, 28'b1111111111111111110101101000, 28'b1111111111111110010110011100, 28'b1111111111111111111000001010, 28'b0000000000000000010010000110}, 
{28'b0000000000000001000010001011, 28'b0000000000000000001010101001, 28'b1111111111111111001000001100, 28'b0000000000000000000000000000, 28'b1111111111111110011111110011}, 
{28'b0000000000000000111011001111, 28'b1111111111111111101001110110, 28'b1111111111111111001001100001, 28'b0000000000000000110101000010, 28'b0000000000000000011000010110}, 
{28'b0000000000000000010001010101, 28'b1111111111111111111000001111, 28'b0000000000000001001100001011, 28'b1111111111111110010001101011, 28'b1111111111111111111010100011}, 
{28'b0000000000000000000000000000, 28'b0000000000000000011110001011, 28'b0000000000000001111100100100, 28'b1111111111111101111011010100, 28'b1111111111111101100001111001}, 
{28'b1111111111111111100110110111, 28'b0000000000000000011100000101, 28'b0000000000000000101101010110, 28'b1111111111111110100100101001, 28'b0000000000000010000101101110}, 
{28'b1111111111111111111111111001, 28'b0000000000000000101010001101, 28'b0000000000000001001000010111, 28'b0000000000000000001001101110, 28'b1111111111111101101101100011}, 
{28'b1111111111111111010100101010, 28'b0000000000000001011101010000, 28'b1111111111111111000110110000, 28'b0000000000000000000001011101, 28'b0000000000000001100011010111}, 
{28'b0000000000000000000110101110, 28'b0000000000000001000100000000, 28'b0000000000000000000111100100, 28'b1111111111111101000000100001, 28'b0000000000000010001100010110}, 
{28'b1111111111111110001010010100, 28'b1111111111111111000001101001, 28'b0000000000000000110110110100, 28'b0000000000000000111110100110, 28'b0000000000000000110011101001}, 
{28'b0000000000000000000001000010, 28'b0000000000000000111101101101, 28'b1111111111111111110110101001, 28'b1111111111111111011001011110, 28'b0000000000000000001000000110}, 
{28'b1111111111111111100101010100, 28'b0000000000000000111111000001, 28'b1111111111111101111111000000, 28'b0000000000000000100011100001, 28'b1111111111111111010111011101}, 
{28'b1111111111111111111011010011, 28'b0000000000000000100100001000, 28'b1111111111111111010100110011, 28'b1111111111111110011001011111, 28'b0000000000000010010111111100}, 
{28'b0000000000000001110010111010, 28'b0000000000000000010001111001, 28'b0000000000000001010011000100, 28'b1111111111111101101001000000, 28'b1111111111111110101111010100}, 
{28'b1111111111111111110000110110, 28'b1111111111111110011101001001, 28'b0000000000000001011101101001, 28'b0000000000000000010010001000, 28'b0000000000000000100000101001}
};

localparam logic signed [27:0] bias [5] = '{
28'b1111111111111111110000000100,  // -0.06223141402006149
28'b1111111111111111101111111100,  // -0.06270556896924973
28'b1111111111111111101110000010,  // -0.07014333456754684
28'b0000000000000000010101000000,  // 0.0820775106549263
28'b0000000000000000110111001011   // 0.2155742198228836
};
endpackage