// Width: 16
// NFRAC: 8
package dense_4_16_8;

localparam logic signed [15:0] weights [32][5] = '{ 
{16'b1111111111111100, 16'b0000000001010000, 16'b1111111110110011, 16'b0000000000010000, 16'b1111111111100100}, 
{16'b1111111101110001, 16'b1111111111110001, 16'b0000000001110101, 16'b1111111111111100, 16'b0000000000000100}, 
{16'b0000000001011111, 16'b0000000000110110, 16'b1111111111111000, 16'b1111111110011000, 16'b1111111111001010}, 
{16'b1111111110011111, 16'b1111111110100000, 16'b1111111111100011, 16'b0000000001001110, 16'b0000000000111100}, 
{16'b0000000000011111, 16'b0000000000100000, 16'b0000000000101000, 16'b1111111111111011, 16'b1111111011111100}, 
{16'b0000000001010011, 16'b1111111110011011, 16'b0000000000101110, 16'b1111111111010110, 16'b1111111111010100}, 
{16'b1111111110011001, 16'b0000000000001001, 16'b1111111111111111, 16'b0000000000101100, 16'b0000000000010001}, 
{16'b1111111111111111, 16'b0000000001001000, 16'b1111111110011011, 16'b0000000000101001, 16'b0000000000100010}, 
{16'b0000000000101001, 16'b1111111111010100, 16'b0000000000000000, 16'b1111111110001001, 16'b1111111111000000}, 
{16'b1111111111111111, 16'b1111111110111011, 16'b0000000000101101, 16'b0000000001101110, 16'b0000000000000000}, 
{16'b1111111111011110, 16'b1111111111011010, 16'b0000000000000000, 16'b0000000010010100, 16'b1111111110111011}, 
{16'b0000000000101011, 16'b0000000000111010, 16'b1111111110101000, 16'b1111111111111000, 16'b0000000000011111}, 
{16'b0000000000000000, 16'b0000000000101010, 16'b0000000000000010, 16'b1111111111001010, 16'b1111111101100000}, 
{16'b0000000000101101, 16'b0000000000010000, 16'b0000000001101011, 16'b1111111111101110, 16'b1111111110010010}, 
{16'b0000000000010111, 16'b1111111111110011, 16'b1111111110100011, 16'b1111111111110111, 16'b0000000010001001}, 
{16'b1111111110000110, 16'b1111111111000001, 16'b1111111111000111, 16'b0000000001100110, 16'b0000000000001000}, 
{16'b0000000001011000, 16'b1111111111010100, 16'b1111111111011101, 16'b1111111111000110, 16'b1111111111110000}, 
{16'b0000000000110001, 16'b1111111111110101, 16'b1111111110010110, 16'b1111111111111000, 16'b0000000000010010}, 
{16'b0000000001000010, 16'b0000000000001010, 16'b1111111111001000, 16'b0000000000000000, 16'b1111111110011111}, 
{16'b0000000000111011, 16'b1111111111101001, 16'b1111111111001001, 16'b0000000000110101, 16'b0000000000011000}, 
{16'b0000000000010001, 16'b1111111111111000, 16'b0000000001001100, 16'b1111111110010001, 16'b1111111111111010}, 
{16'b0000000000000000, 16'b0000000000011110, 16'b0000000001111100, 16'b1111111101111011, 16'b1111111101100001}, 
{16'b1111111111100110, 16'b0000000000011100, 16'b0000000000101101, 16'b1111111110100100, 16'b0000000010000101}, 
{16'b1111111111111111, 16'b0000000000101010, 16'b0000000001001000, 16'b0000000000001001, 16'b1111111101101101}, 
{16'b1111111111010100, 16'b0000000001011101, 16'b1111111111000110, 16'b0000000000000001, 16'b0000000001100011}, 
{16'b0000000000000110, 16'b0000000001000100, 16'b0000000000000111, 16'b1111111101000000, 16'b0000000010001100}, 
{16'b1111111110001010, 16'b1111111111000001, 16'b0000000000110110, 16'b0000000000111110, 16'b0000000000110011}, 
{16'b0000000000000001, 16'b0000000000111101, 16'b1111111111110110, 16'b1111111111011001, 16'b0000000000001000}, 
{16'b1111111111100101, 16'b0000000000111111, 16'b1111111101111111, 16'b0000000000100011, 16'b1111111111010111}, 
{16'b1111111111111011, 16'b0000000000100100, 16'b1111111111010100, 16'b1111111110011001, 16'b0000000010010111}, 
{16'b0000000001110010, 16'b0000000000010001, 16'b0000000001010011, 16'b1111111101101001, 16'b1111111110101111}, 
{16'b1111111111110000, 16'b1111111110011101, 16'b0000000001011101, 16'b0000000000010010, 16'b0000000000100000}
};

localparam logic signed [15:0] bias [5] = '{
16'b1111111111110000,  // -0.06223141402006149
16'b1111111111101111,  // -0.06270556896924973
16'b1111111111101110,  // -0.07014333456754684
16'b0000000000010101,  // 0.0820775106549263
16'b0000000000110111   // 0.2155742198228836
};
endpackage