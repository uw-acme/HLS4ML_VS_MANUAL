// Package with weights and biases for pre-sigmoid dense latency layer
`ifndef SOFTMAX_EXP_PKG
    `define SOFTMAX_EXP_PKG softmax_exp_16_10
`endif
`ifndef SOFTMAX_INVERT_PKG
    `define SOFTMAX_INVERT_PKG softmax_invert_16_10
`endif