// Width: 20
// NFRAC: 10
package dense_3_20_10;

localparam logic signed [19:0] weights [32][32] = '{ 
{20'b11111111111111001101, 20'b11111111111001000000, 20'b11111111111001100000, 20'b11111111111100111100, 20'b00000000000101011111, 20'b00000000000000101100, 20'b11111111111111110010, 20'b11111111111111111111, 20'b11111111111111111111, 20'b11111111111111111111, 20'b00000000000010000001, 20'b11111111110111100100, 20'b11111111111111000010, 20'b00000000001101100011, 20'b11111111111100001000, 20'b11111111110001000100, 20'b11111111111111011010, 20'b00000000000001110010, 20'b00000000000110111101, 20'b11111111111010011011, 20'b11111111101110111100, 20'b11111111111111010000, 20'b00000000000000110010, 20'b11111111111001100011, 20'b00000000000000000000, 20'b00000000010000001100, 20'b11111111101000101100, 20'b11111111111100011101, 20'b11111111111001110010, 20'b11111111111101100110, 20'b00000000000110110001, 20'b11111111111101011100}, 
{20'b00000000001011111101, 20'b00000000011011101011, 20'b00000000000110011011, 20'b11111111110101011110, 20'b00000000000011111010, 20'b11111111111011101000, 20'b11111111111110010000, 20'b00000000010001011100, 20'b00000000000000000110, 20'b11111111111111111111, 20'b11111111111111011111, 20'b11111111110110100101, 20'b11111111111100110001, 20'b00000000001000101001, 20'b11111111011110010011, 20'b11111111111000011101, 20'b11111111111111111111, 20'b11111111111111110111, 20'b11111111111111001010, 20'b11111111111101010111, 20'b11111111111011110111, 20'b11111111111011100110, 20'b00000000000000010001, 20'b11111111111111111110, 20'b11111111111111111001, 20'b11111111101110110110, 20'b00000000000000001100, 20'b00000000000111100010, 20'b11111111111110111111, 20'b11111111110100111101, 20'b00000000000000000010, 20'b00000000000000100110}, 
{20'b11111111110000001111, 20'b00000000000010111100, 20'b00000000000000001010, 20'b00000000000101001010, 20'b11111111110101111010, 20'b00000000000000000000, 20'b00000000000000000001, 20'b11111111110010100100, 20'b00000000001000100100, 20'b11111111111011110011, 20'b11111111111011110110, 20'b11111111101000001101, 20'b11111111111011000001, 20'b00000000001000001011, 20'b00000000000100001110, 20'b11111111111111111110, 20'b11111111111110001010, 20'b11111111111111100111, 20'b11111111110010111101, 20'b00000000000000000011, 20'b00000000000001111111, 20'b00000000000001000110, 20'b00000000000011010110, 20'b00000000001110000101, 20'b00000000000000100110, 20'b11111111110011011000, 20'b00000000001100010001, 20'b00000000000000000000, 20'b00000000000010101001, 20'b11111111111111101001, 20'b00000000000000000000, 20'b00000000100100010011}, 
{20'b00000000001101011001, 20'b11111111111111111111, 20'b11111111111100111000, 20'b00000000010100111100, 20'b00000000010011101001, 20'b00000000000000000000, 20'b00000000000001001011, 20'b00000000001101000001, 20'b11111111111001101010, 20'b11111111111111111111, 20'b11111111110010110100, 20'b00000000000001111010, 20'b00000000000100010000, 20'b11111111110100000010, 20'b00000000000001011111, 20'b11111111111101011100, 20'b11111111111111111111, 20'b11111111111010001011, 20'b00000000000000100111, 20'b00000000000000111000, 20'b00000000000000010000, 20'b11111111111110110101, 20'b00000000010011000110, 20'b00000000001010111110, 20'b00000000001010100010, 20'b00000000000111111100, 20'b00000000001010111011, 20'b00000000000000000000, 20'b11111111111110000111, 20'b00000000001110011111, 20'b00000000000111111111, 20'b11111111111101001100}, 
{20'b00000000010000000000, 20'b11111111111110100000, 20'b11111111110100111010, 20'b11111111100111111100, 20'b00000000001111010001, 20'b00000000000000000000, 20'b11111111110010110111, 20'b11111111110110111101, 20'b11111111111110100000, 20'b11111111100110000110, 20'b11111111011100101001, 20'b00000000001111001000, 20'b00000000010101011001, 20'b00000000010000101111, 20'b11111111101101100110, 20'b11111111100111001100, 20'b00000000000000000000, 20'b11111111111011011110, 20'b00000000000110011011, 20'b00000000000100011100, 20'b11111111111001111110, 20'b11111111111111110010, 20'b00000000010111000101, 20'b11111111010100000000, 20'b00000000000010110100, 20'b11111111101010111011, 20'b00000000000010000110, 20'b11111111111000000011, 20'b11111111110110011100, 20'b11111111111111111111, 20'b00000000000010001111, 20'b00000000010010100100}, 
{20'b00000000000001011000, 20'b11111111111110101011, 20'b11111111110110001011, 20'b11111111110111101010, 20'b00000000001011111001, 20'b00000000000000000000, 20'b11111111110111000011, 20'b11111111111011101001, 20'b11111111110010010011, 20'b11111111111101111100, 20'b11111111111111111111, 20'b00000000000101001000, 20'b00000000000000000000, 20'b00000000001011011100, 20'b11111111101111110100, 20'b11111111111011111010, 20'b00000000000010110110, 20'b11111111110110100111, 20'b11111111111001101011, 20'b11111111111111111111, 20'b00000000000000011000, 20'b00000000001001100101, 20'b00000000001110111100, 20'b11111111111111101010, 20'b11111111111111111111, 20'b00000000001100110100, 20'b11111111101110011010, 20'b11111111111111111111, 20'b11111111111000011011, 20'b11111111111110110100, 20'b11111111111111111001, 20'b00000000000000001101}, 
{20'b00000000000010000101, 20'b11111111110101010111, 20'b00000000000011011101, 20'b11111111111110110001, 20'b11111111111111110000, 20'b00000000000100110110, 20'b11111111111100100110, 20'b11111111101010010101, 20'b11111111111111111111, 20'b11111111111001010101, 20'b11111111110001011000, 20'b00000000001111000111, 20'b00000000000000001110, 20'b00000000010101111001, 20'b00000000011010100001, 20'b00000000000000000101, 20'b11111111111111111111, 20'b11111111110101111010, 20'b11111111111110000001, 20'b00000000001000101111, 20'b11111111100111111111, 20'b00000000000100111111, 20'b00000000001010011100, 20'b00000000000000100110, 20'b00000000000100110011, 20'b00000000100111110010, 20'b11111111110011011000, 20'b11111111111101000110, 20'b11111111111001111011, 20'b00000000001111100101, 20'b11111111111110011011, 20'b11111111111010100101}, 
{20'b11111111101100111010, 20'b00000000000000110000, 20'b11111111101011110111, 20'b00000000001101111011, 20'b00000000100000111001, 20'b00000000000011101101, 20'b00000000000000000111, 20'b00000000000001100000, 20'b11111111111111111111, 20'b00000000000100000110, 20'b00000000101001101000, 20'b11111111111111111111, 20'b00000000001100001100, 20'b00000000010011111011, 20'b00000000011000100110, 20'b00000000100001100110, 20'b00000000000000000000, 20'b11111111110000101100, 20'b00000000001010110000, 20'b11111111111111110100, 20'b11111111101011100101, 20'b11111111111000101111, 20'b00000000000000011011, 20'b11111111111101010110, 20'b11111111101111111101, 20'b00000000111100000001, 20'b11111111111000111110, 20'b00000000000000000000, 20'b00000000000000000000, 20'b00000000011100010000, 20'b00000000000010110101, 20'b00000000001100100010}, 
{20'b00000000001101100000, 20'b11111111111111011000, 20'b00000000000000000000, 20'b11111111111110100111, 20'b00000000000010100111, 20'b11111111111110110010, 20'b11111111111111111111, 20'b00000000000101000001, 20'b00000000000110110000, 20'b11111111110111001110, 20'b00000000000100011110, 20'b00000000000101111111, 20'b00000000000000011000, 20'b00000000001010101001, 20'b11111111111000110011, 20'b11111111100110011111, 20'b00000000000000000000, 20'b11111111111111100011, 20'b11111111111111001001, 20'b11111111110000000010, 20'b11111111111111111101, 20'b00000000000000000000, 20'b11111111111001100000, 20'b11111111111111100011, 20'b11111111111100111101, 20'b00000000000100111111, 20'b00000000001011111101, 20'b11111111111100001011, 20'b11111111111110011011, 20'b11111111111110101101, 20'b00000000000000110111, 20'b11111111110011011100}, 
{20'b11111111111010010100, 20'b00000000001100010011, 20'b00000000000000000000, 20'b00000000000000000000, 20'b00000000011001010110, 20'b00000000001010010011, 20'b11111111111111111111, 20'b11111111101110001111, 20'b00000000000011110001, 20'b11111111101001101011, 20'b11111111010011000110, 20'b11111111111111111111, 20'b00000000000000000000, 20'b00000000001101101110, 20'b00000000000011100011, 20'b00000000000000000000, 20'b11111111110101011111, 20'b00000000000000000000, 20'b00000000000000001101, 20'b00000000000001111100, 20'b00000000000111110011, 20'b11111111111111001011, 20'b11111111110100011110, 20'b00000000000000010000, 20'b11111111111111101000, 20'b00000000100010100110, 20'b00000000001010011100, 20'b11111111111111111111, 20'b11111111111101101110, 20'b00000000010101011000, 20'b11111111111110101110, 20'b11111111111101001100}, 
{20'b11111111101111010000, 20'b00000000000101100110, 20'b11111111111110111000, 20'b11111111111111111111, 20'b11111111111000000111, 20'b11111111110011111010, 20'b00000000000001100010, 20'b00000000000100100111, 20'b11111111111111111111, 20'b11111111111010100001, 20'b11111111101101101011, 20'b00000000000110011011, 20'b00000000001001101110, 20'b00000000000000000000, 20'b00000000011010110110, 20'b11111111101110000001, 20'b00000000000011010100, 20'b11111111110011011111, 20'b00000000001001000001, 20'b11111111111111111111, 20'b11111111111110110001, 20'b00000000000010001111, 20'b00000000000011111011, 20'b00000000000000000000, 20'b11111111110000001100, 20'b00000000000000111111, 20'b11111111101110000111, 20'b11111111111110101110, 20'b11111111111111111111, 20'b00000000010101100111, 20'b11111111111001111010, 20'b00000000000000000000}, 
{20'b11111111111111111111, 20'b00000000000011101011, 20'b00000000000000000000, 20'b00000000001100100001, 20'b11111111111100010000, 20'b11111111111110100111, 20'b00000000000001110111, 20'b11111111111111110100, 20'b11111111111110100001, 20'b00000000010100100000, 20'b00000000010110010111, 20'b00000000000000000001, 20'b11111111110101010110, 20'b11111111101001100001, 20'b11111111111110011000, 20'b00000000000000000000, 20'b00000000000000000000, 20'b11111111111101111101, 20'b11111111110000110000, 20'b00000000001100001111, 20'b00000000000000000100, 20'b00000000001011110111, 20'b11111111111111111111, 20'b00000000010001111111, 20'b00000000000011111101, 20'b00000000001001110011, 20'b00000000001110100100, 20'b11111111111110010110, 20'b11111111110011011110, 20'b11111111110001111001, 20'b11111111111111110101, 20'b11111111101010100110}, 
{20'b11111111111000110000, 20'b11111111111111111111, 20'b00000000000011110100, 20'b11111111110010100110, 20'b00000000000010110000, 20'b11111111111111111111, 20'b11111111111001000011, 20'b11111111111111101100, 20'b11111111111011111111, 20'b00000000000001001100, 20'b00000000000010011111, 20'b11111111111101101101, 20'b00000000000000100001, 20'b00000000000110000000, 20'b11111111101011111111, 20'b11111111111000001010, 20'b00000000000111010011, 20'b11111111111010010101, 20'b00000000000000000000, 20'b11111111111111001100, 20'b00000000000110001011, 20'b00000000000000010000, 20'b11111111111111000000, 20'b00000000000001010111, 20'b00000000001000100111, 20'b11111111111100101011, 20'b00000000000000000000, 20'b11111111110001100010, 20'b11111111111001101111, 20'b11111111111111110001, 20'b00000000000101100011, 20'b00000000000000000000}, 
{20'b11111111101111010111, 20'b00000000001101011100, 20'b11111111111111111111, 20'b11111111111111110010, 20'b11111111111111101100, 20'b00000000000101100111, 20'b11111111111111111111, 20'b00000000011000101101, 20'b11111111111111100001, 20'b11111111111111111111, 20'b00000000000110100101, 20'b00000000000001010011, 20'b00000000000000001101, 20'b00000000000000000000, 20'b00000000000011111001, 20'b00000000001010100100, 20'b00000000000101101100, 20'b00000000000101010101, 20'b11111111111111101110, 20'b00000000001001110101, 20'b00000000000011001110, 20'b00000000000001010010, 20'b11111111111111101110, 20'b00000000001000001000, 20'b11111111111100110100, 20'b11111111110101001001, 20'b11111111111101000010, 20'b11111111111111111111, 20'b00000000000011010000, 20'b00000000000000111100, 20'b00000000000110010000, 20'b00000000001111010101}, 
{20'b11111111111111011001, 20'b11111111110011100010, 20'b00000000000001101001, 20'b11111111111111111110, 20'b00000000011101010100, 20'b11111111111001010111, 20'b11111111101101101101, 20'b00000000000000000000, 20'b00000000000000000000, 20'b11111111111111001011, 20'b00000000000001100011, 20'b00000000001101111110, 20'b00000000001010010011, 20'b00000000000000010101, 20'b00000000000001000100, 20'b11111111111010011010, 20'b00000000000001000100, 20'b11111111111110110010, 20'b00000000000000000000, 20'b00000000000010011010, 20'b11111111111110110011, 20'b00000000000000100111, 20'b00000000001000100001, 20'b00000000000001001011, 20'b11111111111111100111, 20'b11111111110010110010, 20'b00000000000110100000, 20'b11111111111111111111, 20'b11111111111111111111, 20'b11111111111100100110, 20'b11111111111111010100, 20'b11111111111101111111}, 
{20'b00000000000000001110, 20'b11111111111101111110, 20'b11111111111011111101, 20'b11111111111001000000, 20'b11111111101110100000, 20'b00000000010011100000, 20'b00000000000000000000, 20'b00000000000101011001, 20'b00000000001001001011, 20'b00000000000000011010, 20'b11111111111110111010, 20'b00000000001111001110, 20'b00000000000111001010, 20'b11111111110100010011, 20'b11111111111010110011, 20'b11111111111110101011, 20'b11111111110011010000, 20'b11111111111111011100, 20'b00000000000000000000, 20'b11111111111111110110, 20'b00000000000100111111, 20'b11111111111011100111, 20'b00000000000000000000, 20'b00000000000010011101, 20'b11111111111111111111, 20'b11111111110101000100, 20'b00000000000101000000, 20'b00000000000000000000, 20'b00000000000001011011, 20'b00000000000000010110, 20'b11111111110101111000, 20'b00000000000000101010}, 
{20'b11111111111001101110, 20'b11111111111010111101, 20'b00000000000010011100, 20'b11111111111100000001, 20'b11111111111101001000, 20'b00000000000011101101, 20'b11111111111111110101, 20'b00000000000001000111, 20'b00000000000100001100, 20'b11111111111111111111, 20'b00000000000011111101, 20'b11111111111011111011, 20'b11111111111111101100, 20'b11111111111111111111, 20'b00000000000011010011, 20'b11111111111111111111, 20'b00000000001111101000, 20'b11111111111111011100, 20'b00000000000111111100, 20'b11111111111010100100, 20'b00000000000101000100, 20'b00000000000010000000, 20'b00000000000010101100, 20'b00000000000001001010, 20'b11111111111101011001, 20'b11111111110111000101, 20'b11111111110111101101, 20'b00000000000011011101, 20'b11111111111101010100, 20'b00000000000000000001, 20'b11111111111111000111, 20'b00000000000111011011}, 
{20'b11111111111111111111, 20'b11111111110011000010, 20'b11111111110011010011, 20'b11111111111111111111, 20'b00000000010100001100, 20'b11111111111101000110, 20'b00000000000000000000, 20'b00000000001111011101, 20'b11111111111011010001, 20'b00000000000000000000, 20'b11111111110010101000, 20'b11111111110000010100, 20'b00000000001110010110, 20'b00000000000100110101, 20'b11111111111100000111, 20'b11111111110111001111, 20'b00000000000101100001, 20'b00000000000000000000, 20'b11111111111000011001, 20'b00000000000000110110, 20'b00000000000010001110, 20'b11111111111101001010, 20'b00000000001001000101, 20'b11111111100000101001, 20'b00000000000001010011, 20'b00000000000111101001, 20'b11111111111110101011, 20'b00000000000000011110, 20'b11111111111000100010, 20'b11111111111111111111, 20'b11111111111001100100, 20'b11111111111111001110}, 
{20'b00000000000110110011, 20'b00000000001011000010, 20'b00000000010001100111, 20'b11111111111001011101, 20'b00000000001101010100, 20'b00000000001001110011, 20'b00000000000000000001, 20'b00000000001110100100, 20'b00000000001011011011, 20'b11111111111100100101, 20'b00000000010110011100, 20'b11111111110100110100, 20'b00000000010011111000, 20'b00000000001110010010, 20'b11111111011101101010, 20'b11111111111111111110, 20'b00000000000000000000, 20'b00000000000000001011, 20'b00000000001000010100, 20'b11111111101111111001, 20'b00000000000111000101, 20'b11111111111001001101, 20'b11111111110000010011, 20'b11111111111010111110, 20'b00000000001010100010, 20'b11111111101010111000, 20'b11111111110101011100, 20'b11111111111110101011, 20'b11111111111111111111, 20'b11111111101101111100, 20'b00000000001100101001, 20'b00000000000000000000}, 
{20'b11111111111110011011, 20'b00000000000000000001, 20'b11111111111111111111, 20'b11111111111111111111, 20'b11111111110100110000, 20'b00000000000000010010, 20'b00000000000000010000, 20'b11111111111111100001, 20'b11111111111111001110, 20'b11111111111110100001, 20'b00000000000100011100, 20'b11111111111111111110, 20'b00000000000010101001, 20'b11111111110101000011, 20'b00000000000011011010, 20'b11111111111111111110, 20'b00000000000100100000, 20'b00000000001110010100, 20'b11111111110100101101, 20'b00000000000001101010, 20'b11111111111100110101, 20'b00000000000100000111, 20'b00000000000110000101, 20'b11111111111101010001, 20'b11111111110111111101, 20'b00000000000000101010, 20'b00000000011010100010, 20'b11111111111111001110, 20'b11111111111111100000, 20'b00000000001010011000, 20'b00000000000000000000, 20'b00000000011011100101}, 
{20'b11111111101111010011, 20'b00000000000001001010, 20'b11111111111001000100, 20'b00000000001100010000, 20'b00000000000011100000, 20'b11111111111110111111, 20'b11111111111111111111, 20'b11111111111111111111, 20'b11111111110110010011, 20'b11111111111110111100, 20'b00000000000000000000, 20'b11111111101110001110, 20'b00000000000000011001, 20'b11111111111110101110, 20'b11111111111111111010, 20'b11111111111111111111, 20'b11111111111100010001, 20'b00000000000000001011, 20'b00000000000000000110, 20'b00000000000101000100, 20'b00000000000000100011, 20'b00000000000000000000, 20'b00000000000000000000, 20'b11111111111111101111, 20'b00000000000000000000, 20'b00000000000000100101, 20'b00000000010010100110, 20'b11111111111111111111, 20'b11111111111111111111, 20'b11111111111110101100, 20'b00000000000101100110, 20'b11111111111111001011}, 
{20'b11111111111111111100, 20'b11111111111011001010, 20'b00000000000110100010, 20'b00000000000001010001, 20'b11111111110100000110, 20'b00000000000000000001, 20'b00000000001001001001, 20'b11111111111111111111, 20'b00000000000000000000, 20'b11111111111100110110, 20'b00000000000011101011, 20'b00000000000000100110, 20'b00000000001010010110, 20'b11111111101110011101, 20'b11111111111100111110, 20'b11111111111111011100, 20'b00000000000110111010, 20'b11111111110011101101, 20'b00000000000000101011, 20'b11111111100111110110, 20'b11111111111111011001, 20'b11111111111100001100, 20'b11111111111110101101, 20'b00000000001001011101, 20'b11111111111101100111, 20'b11111111110111000000, 20'b00000000000010111001, 20'b00000000000000000000, 20'b00000000001100101010, 20'b00000000010000101111, 20'b11111111110101100000, 20'b11111111110001101000}, 
{20'b00000000000010001010, 20'b00000000000000110100, 20'b11111111110010101111, 20'b11111111111110001011, 20'b11111111111111111111, 20'b00000000000000000100, 20'b00000000000011011001, 20'b00000000001101001010, 20'b00000000000000000000, 20'b00000000000000101001, 20'b00000000000010001111, 20'b11111111101110101111, 20'b11111111111101110111, 20'b11111111101100101011, 20'b00000000001111011000, 20'b00000000000000000000, 20'b11111111111111111110, 20'b11111111101011011111, 20'b11111111111111111111, 20'b11111111111101100111, 20'b11111111111111010101, 20'b00000000000000000000, 20'b00000000000001111111, 20'b11111111111011001100, 20'b00000000000001101100, 20'b00000000001101001001, 20'b00000000001101101001, 20'b00000000001100011111, 20'b00000000001001110110, 20'b00000000000000000000, 20'b00000000000011101001, 20'b00000000011001000100}, 
{20'b11111111111111001100, 20'b11111111111000011000, 20'b00000000001100011101, 20'b11111111111100101101, 20'b00000000000010001110, 20'b00000000000101010111, 20'b11111111111111111111, 20'b11111111110110110100, 20'b11111111111101010001, 20'b11111111101100110001, 20'b00000000001110010100, 20'b00000000000000000111, 20'b00000000001101011010, 20'b00000000010101011100, 20'b11111111111100010001, 20'b11111111100100001000, 20'b11111111111100101011, 20'b00000000001111000010, 20'b11111111110110111100, 20'b11111111111001010100, 20'b00000000000001111001, 20'b00000000000000000010, 20'b11111111101110100011, 20'b11111111111001111000, 20'b11111111111110101111, 20'b11111111111100000110, 20'b00000000000011100101, 20'b00000000010110100000, 20'b00000000000111110110, 20'b11111111111111111111, 20'b00000000000010100101, 20'b00000000000000111000}, 
{20'b00000000000001010110, 20'b00000000001110100001, 20'b00000000000000000000, 20'b00000000001001011101, 20'b00000000011010100110, 20'b11111111111010100010, 20'b11111111111111111111, 20'b11111111111110100101, 20'b00000000001001011000, 20'b11111111111001110111, 20'b11111111111111111101, 20'b00000000001010101010, 20'b00000000000000010001, 20'b00000000000000111000, 20'b11111111001111001000, 20'b11111111111101011101, 20'b00000000000000000000, 20'b00000000000110011011, 20'b11111111111111111001, 20'b00000000001001100011, 20'b11111111111111111111, 20'b11111111111010011110, 20'b11111111101110000001, 20'b00000000000100001011, 20'b00000000001001001001, 20'b11111111011100100000, 20'b11111111111111111111, 20'b00000000000000000000, 20'b00000000010001011010, 20'b11111111100110010110, 20'b00000000000000000011, 20'b11111111111111110011}, 
{20'b00000000000000010011, 20'b11111111110101001000, 20'b00000000000001101110, 20'b11111111111111100001, 20'b00000000000001101010, 20'b00000000010000111011, 20'b11111111101000110011, 20'b00000000000001000110, 20'b00000000001101100011, 20'b11111111110101001101, 20'b11111111111111010000, 20'b00000000000001100100, 20'b11111111111111101101, 20'b00000000000101101110, 20'b00000000000011011011, 20'b11111111111111011101, 20'b00000000000010001001, 20'b00000000000000000000, 20'b00000000000000101100, 20'b00000000001100001001, 20'b11111111111111000110, 20'b11111111110000100000, 20'b11111111101100101001, 20'b11111111111001110011, 20'b11111111101101000110, 20'b00000000000110101010, 20'b00000000010011111100, 20'b00000000001011110011, 20'b11111111111111101010, 20'b11111111110100000100, 20'b11111111110110000011, 20'b00000000000001111010}, 
{20'b00000000000001101010, 20'b11111111110000101101, 20'b11111111111111011101, 20'b00000000000100110100, 20'b11111111110000101100, 20'b00000000000101011011, 20'b11111111111111111111, 20'b11111111111111111111, 20'b11111111111111111111, 20'b00000000000000000000, 20'b00000000001000011101, 20'b11111111111111011100, 20'b00000000000000010011, 20'b00000000000000000000, 20'b00000000000100000100, 20'b11111111111111011101, 20'b00000000000000000101, 20'b11111111111111111110, 20'b11111111110101101100, 20'b11111111101111110100, 20'b11111111111111111110, 20'b11111111101110111010, 20'b11111111110110010111, 20'b11111111110100000110, 20'b00000000011100011111, 20'b00000000000000100100, 20'b11111111111110100001, 20'b00000000001010001001, 20'b00000000011100101110, 20'b00000000001100101000, 20'b11111111011110000100, 20'b11111111111010000100}, 
{20'b00000000001100000001, 20'b11111111111111111111, 20'b00000000001000000010, 20'b11111111111111010111, 20'b00000000001111011110, 20'b11111111111011011011, 20'b00000000000010010001, 20'b00000000001101011000, 20'b00000000001000100100, 20'b11111111101111010010, 20'b11111111111110000001, 20'b00000000000011111011, 20'b00000000000010001101, 20'b11111111111111100010, 20'b00000000000010101101, 20'b00000000000000000000, 20'b00000000001011100110, 20'b00000000000001000111, 20'b00000000001011111110, 20'b11111111111101111001, 20'b11111111111011111011, 20'b11111111111101100110, 20'b11111111111111111111, 20'b00000000001001101010, 20'b11111111111001100001, 20'b11111111111111110011, 20'b00000000000000000000, 20'b00000000000000000000, 20'b00000000000000000000, 20'b00000000001001010110, 20'b11111111110101101111, 20'b11111111111111010000}, 
{20'b11111111111111111110, 20'b11111111111111000000, 20'b11111111110001000111, 20'b00000000001001000110, 20'b00000000000111001001, 20'b11111111111100011111, 20'b11111111111111111111, 20'b11111111111000101111, 20'b00000000000000001101, 20'b11111111111111111111, 20'b11111111110110010110, 20'b11111111111000000111, 20'b00000000001111010101, 20'b00000000000000000000, 20'b11111111111011111010, 20'b11111111111111111111, 20'b00000000000110110110, 20'b11111111111111111111, 20'b11111111111111111111, 20'b11111111111001000101, 20'b00000000001010000111, 20'b00000000000000000000, 20'b00000000000100111111, 20'b11111111111111000101, 20'b00000000000101000001, 20'b00000000000000000100, 20'b00000000000000000000, 20'b00000000000111101101, 20'b11111111111001110110, 20'b11111111111110100001, 20'b00000000000101001000, 20'b11111111111100100111}, 
{20'b11111111111111011101, 20'b11111111110110001000, 20'b00000000010011000001, 20'b11111111111101111010, 20'b00000000000110010010, 20'b11111111110110110110, 20'b00000000000000000000, 20'b00000000000001000110, 20'b11111111110000101010, 20'b11111111111111100101, 20'b11111111111100000010, 20'b00000000000001110111, 20'b11111111110101100000, 20'b00000000000100011010, 20'b00000000000110011110, 20'b00000000000011100000, 20'b00000000000010101111, 20'b11111111111110110010, 20'b11111111101001010101, 20'b11111111111111100100, 20'b11111111111110001011, 20'b00000000000100011110, 20'b11111111111100011100, 20'b11111111111111111111, 20'b00000000000110010100, 20'b11111111111110100010, 20'b11111111111111100010, 20'b00000000001100011100, 20'b11111111110011010000, 20'b11111111110110100011, 20'b00000000001011001110, 20'b00000000000001001001}, 
{20'b00000000001101110010, 20'b00000000000110011100, 20'b00000000000000000001, 20'b11111111111010111010, 20'b11111111111101011111, 20'b11111111111111111110, 20'b00000000000000000000, 20'b11111111111101110010, 20'b11111111111100000001, 20'b11111111111100001101, 20'b00000000000000000000, 20'b00000000000101000100, 20'b00000000000000001101, 20'b00000000000001101100, 20'b11111111111110100100, 20'b00000000000000001011, 20'b11111111111011000101, 20'b00000000000000000001, 20'b11111111111111011011, 20'b11111111111111111110, 20'b00000000000000000100, 20'b00000000000001111001, 20'b00000000000011000111, 20'b00000000000000000000, 20'b00000000000000000000, 20'b11111111101100011101, 20'b11111111111001100111, 20'b00000000000000001101, 20'b00000000000000101001, 20'b00000000000000000010, 20'b11111111111010010101, 20'b00000000000000101011}, 
{20'b00000000000110000000, 20'b11111111011110100100, 20'b11111111111111111111, 20'b11111111111101100101, 20'b11111111111000100011, 20'b11111111111111101100, 20'b00000000000000000000, 20'b00000000010001100001, 20'b11111111111110100110, 20'b11111111111111010011, 20'b00000000000010101000, 20'b11111111101010110110, 20'b00000000000000110001, 20'b11111111110001111110, 20'b00000000010111000111, 20'b11111111111110010100, 20'b11111111111000110000, 20'b11111111101110011111, 20'b11111111111111101010, 20'b11111111101001010110, 20'b11111111100110000101, 20'b11111111111111111111, 20'b00000000000000000000, 20'b00000000000000000000, 20'b00000000000111110011, 20'b11111111111111100011, 20'b11111111110110011101, 20'b11111111111101101011, 20'b11111111111111010000, 20'b00000000000000000000, 20'b11111111111110111111, 20'b11111111101001100110}
};

localparam logic signed [19:0] bias [32] = '{
20'b00000000001000011100,  // 0.5280959606170654
20'b00000000001101011101,  // 0.8414360880851746
20'b00000000000110010111,  // 0.397830605506897
20'b00000000000110100100,  // 0.4105983078479767
20'b11111111000101011110,  // -3.657735586166382
20'b11111111110001101000,  // -0.8977976441383362
20'b00000000011011010010,  // 1.7051936388015747
20'b11111111101011100100,  // -1.2765135765075684
20'b11111111110110101010,  // -0.5837795734405518
20'b00000000101011001100,  // 2.699671983718872
20'b00000000000011011110,  // 0.2170683741569519
20'b00000000001110000110,  // 0.8814588785171509
20'b11111111010101110110,  // -2.634300947189331
20'b11111111100001111101,  // -1.877297282218933
20'b00000000011010100110,  // 1.6625694036483765
20'b00000000101011111011,  // 2.7459704875946045
20'b11111111111000010110,  // -0.47838035225868225
20'b00000000011011001011,  // 1.6984987258911133
20'b00000000001101101011,  // 0.8548859357833862
20'b00000000010000000100,  // 1.0045719146728516
20'b00000000010110101101,  // 1.4197649955749512
20'b00000000001101010100,  // 0.832463800907135
20'b00000000001000101100,  // 0.5434179306030273
20'b00000000001110110101,  // 0.9277304410934448
20'b11111111111010100001,  // -0.3426123857498169
20'b11111111110111000011,  // -0.5587119460105896
20'b11111111110110000100,  // -0.6208624839782715
20'b11111111101011100001,  // -1.2802538871765137
20'b00000000000000111100,  // 0.05940237268805504
20'b11111111110010110110,  // -0.8213341236114502
20'b00000000001110000011,  // 0.8783953189849854
20'b11111111110000110011   // -0.949700653553009
};
endpackage