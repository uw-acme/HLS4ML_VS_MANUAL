//Width: 37
//Int: 13
package dense_1_gen;

localparam logic signed [36:0] weights [16][64] = '{
{37'b0000000000000010000010100101000111100, 37'b1111111111111010110010010011011110110, 37'b1111111111111110100011011110010010000, 37'b1111111111111110001100000011010000000, 37'b1111111111111100110000101000011111111, 37'b0000000000000000111000100000001101110, 37'b1111111111110111101101000011101011100, 37'b0000000000000000000000000011111100001, 37'b0000000000000000011101101111011011100, 37'b0000000000000010000110111011111000100, 37'b0000000000000000000001100000110000111, 37'b1111111111111100110000110111101111111, 37'b1111111111111111111111011100110111101, 37'b0000000000000001101011000011001100011, 37'b0000000000000000010001001001110111001, 37'b1111111111111101111010000011000101001, 37'b0000000000000001110111001100011010110, 37'b0000000000000000011110000010000010000, 37'b0000000000000000000000000010011000010, 37'b1111111111111111111111111011011000010, 37'b0000000000000011000000111111101100100, 37'b1111111111111101010110010011011000110, 37'b1111111111111111110100101101101010010, 37'b0000000000000011110010000001010100010, 37'b1111111111111101011011011001110000101, 37'b1111111111111010100010100000001010010, 37'b1111111111111101110010111110100100111, 37'b1111111111111110011100000010111010111, 37'b1111111111111111001010011101001001100, 37'b1111111111111111111111000110101001010, 37'b0000000000000000010011010100001010110, 37'b0000000000000001111101101001011000010, 37'b0000000000000001100100001110101011010, 37'b1111111111111111111001010010110100111, 37'b0000000000000000000000000100110011010, 37'b0000000000000010011111011100101000010, 37'b1111111111111111110110110001111010011, 37'b1111111111111101111111011000100010000, 37'b0000000000000000001101111101001101000, 37'b0000000000000001100010100101011100100, 37'b1111111111111111111001110110111101100, 37'b0000000000000010001100111000101011100, 37'b1111111111111101110111100110001011111, 37'b0000000000000111011011100001001110000, 37'b1111111111111111111111011100111100011, 37'b0000000000000011100111101101101011010, 37'b0000000000000000000000000001110100100, 37'b0000000000000001011110011001100000101, 37'b0000000000000001100100011001110111010, 37'b1111111111111111110011111111100101101, 37'b0000000000000000000000000001111100111, 37'b0000000000000001010010001001001000111, 37'b0000000000000001101110100011111101011, 37'b0000000000000000100111110100000100110, 37'b1111111111111111000100111111101100111, 37'b1111111111111101100001000110100001100, 37'b0000000000000100010010101000000101000, 37'b1111111111111100000000001101011101111, 37'b0000000000000011101111011100001100110, 37'b1111111111111101001010100100111101011, 37'b0000000000000110010110000101001010100, 37'b1111111111111111111100001110000111101, 37'b0000000000000000000101110111011000001, 37'b0000000000000000101001100010100110001},
{37'b0000000000000000000001011100011100111, 37'b1111111111111101011011110000011011011, 37'b1111111111111110111100001100001000100, 37'b1111111111111101110000110111010100101, 37'b1111111111111101011101011110111011000, 37'b0000000000000000110110100111111011100, 37'b1111111111111001111101101110010001110, 37'b1111111111111111111110110110110000000, 37'b1111111111111110001011101000011111011, 37'b0000000000000001011000010000111110110, 37'b0000000000000000000011011000011100001, 37'b1111111111111111010011111000100101011, 37'b0000000000000001100100111011011001100, 37'b0000000000000000000000000010000101101, 37'b1111111111111111111111111011010110000, 37'b0000000000000001101010010011011000000, 37'b1111111111111111111100111011010000111, 37'b0000000000000000000000001010111010101, 37'b1111111111111110100010101110011011001, 37'b1111111111111101111111111001011111000, 37'b0000000000000011100010011111100101100, 37'b1111111111111111010110100100011111000, 37'b0000000000000000011000100011000010100, 37'b0000000000000101100101110100110001101, 37'b0000000000000010000011110110110010001, 37'b1111111111111110001010000101010001101, 37'b1111111111111110001001110001101010011, 37'b1111111111111111111111110101001110011, 37'b1111111111111111001100000011101100100, 37'b1111111111111100110000011111100101101, 37'b1111111111111111100001010110011011000, 37'b0000000000000011101000111010001100111, 37'b0000000000000010001110101001001101010, 37'b0000000000000100011001101011111101110, 37'b0000000000000101000010000100010000101, 37'b0000000000000000011001110110011010110, 37'b1111111111111111000011011000100001111, 37'b1111111111111100100001110010001000011, 37'b0000000000000000011101000000011001000, 37'b0000000000000001100000101101100001010, 37'b0000000000000000001011101111100110101, 37'b0000000000000001101001101101001100111, 37'b1111111111111110010011001001100001001, 37'b0000000000000010000001000001001011010, 37'b0000000000000001011000001111100001000, 37'b0000000000000000011001100001001101001, 37'b1111111111111101010001111101010111001, 37'b0000000000000000101000101101100001100, 37'b0000000000000010000101011111000101100, 37'b0000000000000000001111010101111011011, 37'b0000000000000000001100101110001111101, 37'b0000000000001001010000100000111000010, 37'b1111111111111111011001101111010011010, 37'b1111111111111111001101110100010010100, 37'b1111111111111111100100001100010110101, 37'b1111111111111111111100000001011110100, 37'b0000000000000010000011100011001011000, 37'b1111111111111101000010100110101000011, 37'b0000000000000111111000011111100001101, 37'b0000000000000000000010011101010000101, 37'b0000000000000100001010100011001101111, 37'b0000000000000001111010111111001010010, 37'b0000000000000110100101001110011100100, 37'b0000000000000001001000001101011010001},
{37'b1111111111111111111100000110001101011, 37'b0000000000000000000000000000101000100, 37'b1111111111111111010101011011000010101, 37'b1111111111111110100101111001100011011, 37'b1111111111111110100001011111100100001, 37'b0000000000000000010101011011101010110, 37'b0000000000001011110110001111100110010, 37'b1111111111111111111111111110101101011, 37'b1111111111110101110111110010010001100, 37'b1111111111111111111111111100111000100, 37'b1111111111111111111111000111010111001, 37'b1111111111111111110110110101101000010, 37'b1111111111111110001011100101010110100, 37'b0000000000000000000000101001111000101, 37'b1111111111111111111011001100111101001, 37'b0000000000000001010110000100011011000, 37'b0000000000000111001111100101011000000, 37'b1111111111111111111111111110001000000, 37'b0000000000000000100100111111100011000, 37'b0000000000000000000000001010000011010, 37'b0000000000000011010011000010100000000, 37'b1111111111111010001110101111010100110, 37'b0000000000000100100111101011100111101, 37'b1111111111111010010010100101010010111, 37'b0000000000000111100101101000111000100, 37'b1111111111111101001110101000111000110, 37'b1111111111111110000010101010101000011, 37'b1111111111111010010000100111011101100, 37'b0000000000001010001100000011110011100, 37'b0000000000000010001101001110101100010, 37'b0000000000000000000101110101101010011, 37'b0000000000000100001001000100110101000, 37'b0000000000001000001010011100101100100, 37'b1111111111110110011100001011110100000, 37'b1111111111111111001111000100010010010, 37'b0000000000000000010000010110100101001, 37'b1111111111111110001001101111100111111, 37'b0000000000000111001011010001100111110, 37'b1111111111111111101011110110000010001, 37'b0000000000000010100000010011001000000, 37'b0000000000000010101010100010100100110, 37'b0000000000000010111101010010100011011, 37'b1111111111111111111111111110010110111, 37'b1111111111111111111111111010100000011, 37'b1111111111111111110111001010100111011, 37'b0000000000000001010000011100111001110, 37'b1111111111111101110000110000110011111, 37'b1111111111111110101000110100011110010, 37'b1111111111111111110111000100010011000, 37'b0000000000000011001001011000111101100, 37'b1111111111111110100101111011101011001, 37'b0000000000000001001100111000000100101, 37'b1111111111111111111111110001010100010, 37'b0000000000000001000100101111010001000, 37'b1111111111111110100110001001110000001, 37'b1111111111111111111111111100111001010, 37'b1111111111111101100010001000101001000, 37'b1111111111111010101001001101000111101, 37'b1111111111111111111110111110010001101, 37'b0000000000000000000000000001011010001, 37'b0000000000001100010101111100010110110, 37'b0000000000000000000110101010010001000, 37'b1111111111111111111110101000111010010, 37'b1111111111111101100001100100111010001},
{37'b1111111111111100010101011010111001010, 37'b1111111111111101000011010010000000111, 37'b1111111111111010011101010110100100000, 37'b0000000000000010011101110100100110100, 37'b1111111111111101011110010001101100111, 37'b1111111111110101001110101110010011000, 37'b1111111111111111000101010001111000010, 37'b1111111111111101100010010001111111111, 37'b0000000000000001110010101110001011110, 37'b1111111111111111111111111111100011000, 37'b0000000000001010000111111001001001100, 37'b1111111111111111001001111110111011010, 37'b1111111111111001101111011001011001101, 37'b0000000000000100101000100100101011101, 37'b0000000000000000001100111000110000100, 37'b1111111111111111111111001110110111100, 37'b1111111111111100011100110011111001001, 37'b1111111111111111111111111110011011100, 37'b0000000000000000000000000010110001000, 37'b1111111111111110001100001111111110001, 37'b1111111111110110110010101110101010010, 37'b1111111111111111000110110110000010011, 37'b1111111111111010011010011110011011111, 37'b0000000000000001100101100110110111001, 37'b1111111111111100111001111100101100001, 37'b1111111111111000101000101000011101100, 37'b0000000000000010100000001001011001100, 37'b0000000000000101111001001001001000000, 37'b0000000000001010010111001011000111010, 37'b1111111111111100010100100000000111111, 37'b1111111111111011010101101100000011001, 37'b0000000000000000100101110100000010100, 37'b0000000000000100000000000101110000110, 37'b1111111111111001010001010000000101110, 37'b1111111111111101011111000000100010101, 37'b0000000000000000000000000000000001010, 37'b1111111111111010001100010001110100011, 37'b0000000000000001111100001010011100100, 37'b1111111111111100011110001001100110001, 37'b0000000000000000111101000111100101001, 37'b0000000000000011101010110011000101100, 37'b0000000000000001010000010000111011000, 37'b0000000000000000000000000000000000111, 37'b0000000000000000001010011010000101111, 37'b0000000000000100011010111001101100011, 37'b1111111111111110011001101000101011110, 37'b1111111111111111111111111100011111011, 37'b1111111111111101001111111001111111101, 37'b1111111111111111111111111100001111011, 37'b1111111111111111001110011110100100001, 37'b1111111111111011000100111010000010101, 37'b0000000000000000101100011100000000101, 37'b1111111111111111111111111101100011000, 37'b0000000000000001101111101100010101001, 37'b0000000000000010100001011110110010000, 37'b0000000000000101001011010101100010000, 37'b1111111111111000010000100111110101111, 37'b1111111111111000100100011101101100101, 37'b1111111111111010010110111111110000001, 37'b0000000000000110111011100000010011101, 37'b0000000000001101111111100011011101100, 37'b1111111111111000110011011001101101001, 37'b1111111111111111100100010010111101011, 37'b0000000000000011011110010110011100011},
{37'b0000000000000010101111001100100110110, 37'b1111111111111011000011010110000101100, 37'b1111111111111101111011001110001111011, 37'b1111111111111111111111111111100111000, 37'b1111111111111110110001001010000111101, 37'b0000000000000010101110001101101001111, 37'b0000000000000001100001000001100101100, 37'b1111111111111111111111111011100010101, 37'b1111111111111011001110001010001010101, 37'b1111111111111110000100001111110001111, 37'b1111111111111101000011001111010101001, 37'b0000000000000000011011000111000111101, 37'b0000000000000000000000101001011110001, 37'b0000000000000000000000000001001011000, 37'b1111111111111111101011010001101100101, 37'b0000000000000010110111000111111011110, 37'b0000000000000001000100011011001010010, 37'b1111111111111100110110110110011000111, 37'b0000000000000000001111101100100111111, 37'b0000000000000000000110111011001010001, 37'b0000000000000001101011100110101111110, 37'b1111111111111111000011100100101010001, 37'b0000000000000000100110000111000110100, 37'b1111111111111111110110001111100011111, 37'b0000000000001000100001101101011101100, 37'b1111111111111110100000100110100111101, 37'b1111111111111101110000000010110001010, 37'b1111111111111100110001010101001010100, 37'b0000000000000000000000000010000100001, 37'b0000000000000001010100010110010100110, 37'b0000000000000000111011100000110000010, 37'b0000000000000010001100000100000110000, 37'b1111111111111111111001101000101110001, 37'b0000000000000000100101111100111110000, 37'b0000000000000001000010111010101100111, 37'b1111111111111111111111111111010111100, 37'b0000000000000000000011001011101001100, 37'b0000000000000111000011010110111011011, 37'b1111111111111101101100000110111110101, 37'b1111111111111111011000110001001111101, 37'b0000000000000011011101110100001101001, 37'b0000000000000001111111011000101001000, 37'b1111111111111100000101101010011100011, 37'b0000000000000000000011000000100100010, 37'b1111111111110111011101000000101000010, 37'b1111111111111111111111111110011000111, 37'b1111111111111111000001010001000011011, 37'b0000000000000000000110000111101010000, 37'b1111111111111111111111111010001101101, 37'b1111111111111111110011111111110110101, 37'b1111111111111111111111111110100001000, 37'b0000000000000001100000010011000001010, 37'b1111111111111111111101011000001110001, 37'b0000000000000010100010101100010110010, 37'b1111111111111110011110001001100001000, 37'b1111111111111010000111100110010000100, 37'b1111111111111100010001001100100011011, 37'b1111111111111011111011001100100010010, 37'b1111111111111011000101101100111011011, 37'b0000000000000101111110011011101000010, 37'b0000000000001010111111010011111101110, 37'b0000000000000110010101111101101010001, 37'b0000000000000000111110110000011000010, 37'b1111111111111111111111111010101011000},
{37'b1111111111111100011011110111010111011, 37'b1111111111111010111101001000100011010, 37'b0000000000000000000000000100001010010, 37'b0000000000000010011101010010111001001, 37'b0000000000000010010010000100000101010, 37'b1111111111111110010011011011011100111, 37'b0000000000000100101010000101100110000, 37'b1111111111111111111111111100101111111, 37'b0000000000000001111100110000001101100, 37'b1111111111111111111111111110100101100, 37'b1111111111111111111011001101100101011, 37'b1111111111111111011010110100111000110, 37'b1111111111111110100101101011110110000, 37'b0000000000000100101000000001100101101, 37'b1111111111111111010010010011101001010, 37'b0000000000000000000000000110011100010, 37'b1111111111111011000000000101001000011, 37'b1111111111111101001010100011010011011, 37'b0000000000000000000000000100001010100, 37'b1111111111111111111111111100000010001, 37'b1111111111111111100111101001011110111, 37'b1111111111111101011111010100111011010, 37'b1111111111111101011100110010111010101, 37'b0000000000000011101110010011001101000, 37'b1111111111111101011101001010100111101, 37'b1111111111111111111111100011001110111, 37'b0000000000000010000011001000100101000, 37'b1111111111111111011010100110000001010, 37'b1111111111111000100010011011001001100, 37'b1111111111111111111111111101100001101, 37'b1111111111111111011101110001000000101, 37'b1111111111111111111010101111011010000, 37'b1111111111111111111010000100010010011, 37'b0000000000000000010100111100101110010, 37'b0000000000000001000011100010001011010, 37'b0000000000000010110001000000011001000, 37'b0000000000000000000110111101110001101, 37'b1111111111111111001101110010011100110, 37'b1111111111111101111001100011010010010, 37'b1111111111111111111111000010100010100, 37'b1111111111111110101001011100110011011, 37'b1111111111111011110011110011001110010, 37'b0000000000000011001100111110010101000, 37'b0000000000000000000101100000101111000, 37'b0000000000000100110100111011101010110, 37'b0000000000000000000000000000011110001, 37'b1111111111111111111111111011011101110, 37'b0000000000000000110000101011111000010, 37'b1111111111111100101001011001111100101, 37'b0000000000000001110111110100011001110, 37'b0000000000000000000000000000010110011, 37'b1111111111111111001100010000010111110, 37'b1111111111111101000110111110111001111, 37'b0000000000000011000101111001011000110, 37'b1111111111111111111111111111010000011, 37'b0000000000000010110001101100101000010, 37'b0000000000000001101110111010010010001, 37'b0000000000000001101000011001101100111, 37'b1111111111111111110110011101001111111, 37'b1111111111111111111011110001010110000, 37'b1111111111111001100010001010100111000, 37'b1111111111111110111111011000001110000, 37'b1111111111111111100010110001100111100, 37'b1111111111111111111111110011000001001},
{37'b1111111111111101101111001101100101111, 37'b1111111111111101010100011011010010101, 37'b1111111111111100100011000011101001010, 37'b1111111111111111011100011000000100101, 37'b1111111111111110111011110001110011100, 37'b0000000000000000110101011000000010001, 37'b1111111111111010011010100010010110111, 37'b1111111111111110110011001010010100011, 37'b1111111111111110001101001011100100111, 37'b1111111111111111111111111010011001100, 37'b1111111111111101101100110101101100011, 37'b0000000000000010110010001000001110110, 37'b0000000000000000010010001111000100010, 37'b0000000000000001000110100010100111110, 37'b0000000000000010011111101111110010010, 37'b0000000000000000000000001001001010100, 37'b0000000000000110011000001010011101000, 37'b0000000000000000101101110000001111110, 37'b0000000000000001111100010101111110110, 37'b0000000000000010001001011101101110101, 37'b1111111111111110101111110000110001001, 37'b0000000000000010111010000010111010000, 37'b1111111111111110000011110000000101011, 37'b1111111111111011111111000001101110100, 37'b0000000000000001011000110000000101000, 37'b0000000000000100001000100101010101000, 37'b1111111111111111111101110111010100010, 37'b0000000000000000011011100101010010000, 37'b1111111111111000011001001010100010011, 37'b0000000000000010010010101100111111000, 37'b0000000000000010001000110010101110100, 37'b1111111111111101000000111000001101110, 37'b0000000000000011110001011001100010010, 37'b0000000000000101010100010100000010101, 37'b0000000000000000000000000001101111000, 37'b0000000000000010101111010010011011101, 37'b1111111111111111111111111110011011111, 37'b0000000000000010010001100011101101110, 37'b0000000000000001100101111101111101010, 37'b0000000000000000000000000000010000000, 37'b1111111111111111000011101000111001100, 37'b1111111111111101000101110100001001001, 37'b0000000000000001001001011100111111101, 37'b0000000000000011110111011111011100000, 37'b0000000000000100001001110001001111001, 37'b1111111111111110101001111010101011100, 37'b1111111111111111010101010001000000101, 37'b1111111111111110011110110010100111111, 37'b1111111111111110111010110000010001001, 37'b0000000000000000111100100111101011100, 37'b0000000000000000000001101000110000111, 37'b0000000000000000010001011101011000010, 37'b0000000000000000000000000000110010010, 37'b0000000000000001011100110111110000010, 37'b1111111111111110100110101001110101101, 37'b0000000000000110001010101101000101101, 37'b0000000000000010110110010001110110010, 37'b1111111111111111110011010111011111001, 37'b0000000000000011000111110101101010000, 37'b0000000000000001101111001000011001101, 37'b1111111111110010111111111111110101110, 37'b1111111111111011011000111101001100101, 37'b1111111111111110100111110100011110111, 37'b1111111111111111111010111000001010101},
{37'b0000000000000000000010101000101100110, 37'b0000000000000001111010011111011011100, 37'b1111111111111111111111110100110011001, 37'b1111111111111111111111101110111011010, 37'b1111111111111101011011000011111000001, 37'b1111111111111111110000000001110011010, 37'b1111111111111101111100001111111111100, 37'b0000000000000000000000000011111001101, 37'b0000000000000000001110000111101011111, 37'b0000000000000011000111000101011110110, 37'b0000000000000000000111011110110100101, 37'b1111111111111100111110100000100100101, 37'b1111111111111111011111111111011001000, 37'b0000000000000000000000000101011001011, 37'b1111111111111111100101000000100001111, 37'b1111111111111100011001110010111001011, 37'b1111111111111001001101100111101111110, 37'b1111111111111111111111110110111010000, 37'b1111111111111011001010100110101010000, 37'b1111111111111100011011101101110011111, 37'b1111111111111100111000100100010111100, 37'b0000000000000010110001110001000111000, 37'b0000000000000000011000000010000011000, 37'b1111111111111110110111000101001011111, 37'b1111111111111100100000010001010001101, 37'b0000000000000001001111100100100000101, 37'b0000000000000000000000000000110100110, 37'b0000000000000011111111101011111000100, 37'b0000000000000110011100101010100010011, 37'b1111111111111111101011011010101010110, 37'b0000000000000000000000010111101011110, 37'b0000000000000001110110000011111100000, 37'b1111111111111010100010101110001111011, 37'b1111111111111101000010000111000011001, 37'b0000000000000000011100011100000010010, 37'b0000000000000000101111011010010001001, 37'b1111111111111101110000010111110001111, 37'b0000000000000001111010101001000111100, 37'b0000000000000001000011100111011110010, 37'b1111111111111110110001110011111010100, 37'b1111111111111100101001000011010111001, 37'b1111111111111111101101000011001011100, 37'b0000000000000000010000110010111001111, 37'b1111111111111110101010111101000011101, 37'b0000000000000000011100100100010111100, 37'b0000000000000001110101011011010010000, 37'b1111111111111111000010111000100000011, 37'b0000000000000000001100001110110010111, 37'b0000000000000000000000000001011100110, 37'b1111111111111110010000011111100101001, 37'b1111111111111100111001001111101110101, 37'b0000000000000011010100111111111001000, 37'b0000000000000001000000111111101110101, 37'b1111111111111110100100110011110000100, 37'b0000000000000001000011110111110110010, 37'b1111111111111111100000011010001010111, 37'b1111111111111100001101000101010011111, 37'b1111111111111110111011110001011101010, 37'b1111111111111111100101010000011110111, 37'b1111111111111111011100000101111111111, 37'b0000000000000110101001001010111000001, 37'b0000000000000001100001101111010010000, 37'b1111111111111111100111001100101001111, 37'b1111111111111111111111110101010010101},
{37'b0000000000000000000111100001100111110, 37'b0000000000000100101100011110000111010, 37'b1111111111111011010110101101111000000, 37'b1111111111111110001001101101101100001, 37'b0000000000000010100101001100010011010, 37'b1111111111111110010110011110011100110, 37'b0000000000001001101100001000101010010, 37'b1111111111111101101100101101110111011, 37'b1111111111111111111111111011010010101, 37'b0000000000000010010110001001101101010, 37'b0000000000000010000010001011010000110, 37'b1111111111111111111110101110100000000, 37'b1111111111111111100111011010110001000, 37'b1111111111111100001001001010110101101, 37'b0000000000000010010000000100110110110, 37'b0000000000000001010001110010101111010, 37'b1111111111111110011100110001011101011, 37'b1111111111111111111111111111001111000, 37'b0000000000000000000000000000110010001, 37'b0000000000000000000000001001111001110, 37'b0000000000000010000111110111001000010, 37'b1111111111111100010100101001101000101, 37'b0000000000000011001000110011010100000, 37'b0000000000000100111001110001000101001, 37'b1111111111111111010011010101001100101, 37'b1111111111111111111111110111010010100, 37'b1111111111111111110111101010100010000, 37'b1111111111111111111111111001001101101, 37'b0000000000000101111000111011110101100, 37'b0000000000000000000010100010100111111, 37'b1111111111111101110100000111011001010, 37'b0000000000000000000000000000011101000, 37'b0000000000000011000100101101110110100, 37'b1111111111111001100000110001000011010, 37'b1111111111111011101011001011001011011, 37'b0000000000000001100101110000000111011, 37'b0000000000000001000110111010000011000, 37'b1111111111111011011011011010010001011, 37'b1111111111111110011111001001110000101, 37'b1111111111111110010010010100010111011, 37'b0000000000000011001101010101001011001, 37'b0000000000000011001000001010100000101, 37'b0000000000000000000000000011000110100, 37'b1111111111111101110101110001000000001, 37'b0000000000000000000000011010101110000, 37'b0000000000000011001010011100010001110, 37'b1111111111111111100001110101000010101, 37'b1111111111111111111111111011000111101, 37'b0000000000000000000101111000101001001, 37'b0000000000000001111101011101111011100, 37'b1111111111111111100010100110101101001, 37'b1111111111111110011100111000000001010, 37'b0000000000000010110000001110110100010, 37'b1111111111111110010001111010101001101, 37'b0000000000000010001111001101100010000, 37'b0000000000000100101011010110100111000, 37'b0000000000000000010100011111011010000, 37'b0000000000000010000110111101111100111, 37'b1111111111111100110011000110011001001, 37'b1111111111111101000100001000001000101, 37'b0000000000000110101001111011000100110, 37'b1111111111111110111110000100000010110, 37'b0000000000000000010111100001011111110, 37'b1111111111111111010000001000101000101},
{37'b0000000000000000001000010010111110010, 37'b1111111111111100011000010111001001001, 37'b0000000000000010111100110111100110010, 37'b1111111111111101101110101001011001001, 37'b1111111111111111111110011111110001110, 37'b0000000000000001101100010010101001100, 37'b1111111111111011010110000010011101111, 37'b0000000000000001100010000001011011111, 37'b0000000000000011111011001000000100000, 37'b0000000000000001001110111100110011100, 37'b0000000000000010111001100001100100100, 37'b0000000000000010100101001000100101000, 37'b1111111111111101100011111111011010000, 37'b1111111111111111011001001001110110111, 37'b1111111111111111100101101011111111111, 37'b0000000000000000000000100110110011101, 37'b1111111111111000010100101001011101011, 37'b0000000000000010100101011101100101010, 37'b1111111111111111101101011110111000011, 37'b0000000000000000001111111010110110100, 37'b1111111111111101001011100000100110011, 37'b0000000000000000100011110001110010101, 37'b0000000000000001001110011000100101101, 37'b1111111111111111111111110100000101010, 37'b1111111111111100010100010110001001001, 37'b1111111111111111100111100011001111010, 37'b1111111111111111010110000001100110010, 37'b0000000000001001111110111011001110000, 37'b1111111111111010101100110011110111110, 37'b0000000000000000100010000001011001001, 37'b0000000000000000110001101011001001010, 37'b1111111111111111100010000101010001011, 37'b1111111111111110001110111000011100001, 37'b0000000000000000111011101011110001001, 37'b1111111111111111010111111100111011000, 37'b1111111111111110111011001100101111011, 37'b1111111111111110100100110111111110010, 37'b1111111111111110010100011101001101100, 37'b1111111111111111110100101100001111011, 37'b1111111111111101100111101101111001010, 37'b0000000000000010100100110000110101000, 37'b0000000000000000111111001100000100111, 37'b0000000000000011111110010111000011100, 37'b0000000000000000101100111010101100101, 37'b0000000000000000010010111000101001101, 37'b1111111111111101101011000100100110111, 37'b0000000000000000000000000000101011010, 37'b1111111111111111111111111010010001100, 37'b1111111111111111111111110000110111110, 37'b0000000000000001100011001111110000110, 37'b0000000000000001011010110110010100111, 37'b0000000000000010010110111110010011110, 37'b1111111111111111111100111001001001001, 37'b1111111111111101101001110010010110110, 37'b0000000000000000000100100111100001100, 37'b0000000000000000000000000011110000001, 37'b0000000000000010100101000110001111111, 37'b1111111111111110011001001001000001011, 37'b1111111111111011100110001010001110111, 37'b0000000000000100011111011000010000101, 37'b1111111111111101101001100010110111110, 37'b0000000000001001010011111000000101110, 37'b1111111111111111110101110111000110111, 37'b1111111111111101001010100000001000001},
{37'b1111111111111011011000111111111001111, 37'b1111111111111111111111000010101011000, 37'b1111111111111100101110010011000100010, 37'b0000000000000001110101111110111010100, 37'b0000000000000010000110110110010010110, 37'b1111111111111111001011100111111111011, 37'b0000000000000100001000101101111010110, 37'b1111111111111110101000110001010110111, 37'b1111111111111100001010100100011001111, 37'b1111111111111101000100001000100101110, 37'b1111111111111101111111011000111110111, 37'b1111111111111100001100010111001010101, 37'b1111111111111110001010110011100010011, 37'b0000000000000001100100110101110110100, 37'b0000000000000000000000000001110001001, 37'b0000000000000000000000001000101100010, 37'b0000000000000110101111011001001100101, 37'b1111111111111111101001111001000001010, 37'b1111111111111111111111011101010010101, 37'b0000000000000011010010100011011010000, 37'b0000000000000010010101111011110100010, 37'b1111111111111011010111101110000111100, 37'b1111111111111100111100001110110101001, 37'b0000000000000001100000110010010011001, 37'b1111111111111100100011100010000001011, 37'b1111111111111111110101010001001111100, 37'b1111111111111101111011000110011000001, 37'b1111111111111101010100111010101000000, 37'b1111111111111100100000111100100110101, 37'b0000000000000010011010101110010111010, 37'b0000000000000001110100101000010110011, 37'b1111111111111110110000001010101000100, 37'b1111111111111111011010110011100010000, 37'b1111111111111000001101010101101010110, 37'b1111111111111110100101100010101101111, 37'b0000000000000000011001010100011111010, 37'b1111111111111110111101101011101011100, 37'b1111111111111101101000001100100001101, 37'b1111111111111111111110001001110010110, 37'b0000000000000000111100111001110110000, 37'b1111111111111111000011000000111111110, 37'b1111111111111111111110101010111101010, 37'b1111111111111111101110000110010000110, 37'b1111111111111010101011111111011110000, 37'b0000000000000000000000011011100000111, 37'b0000000000000000000000000001101011010, 37'b0000000000000010101110001000010001001, 37'b1111111111111111000000010111100100100, 37'b0000000000000011011000111011101011000, 37'b1111111111111110011110011100001000111, 37'b0000000000000010010011011110011010001, 37'b1111111111111111111111010001011000110, 37'b0000000000000001110011100111110000110, 37'b1111111111111100110111101010111011111, 37'b1111111111111111111111111111000111101, 37'b0000000000000100000110001000110010010, 37'b0000000000000010100000000111110010101, 37'b0000000000000010010101100011111100110, 37'b0000000000000000001100111110000110000, 37'b1111111111111100110011010010000000010, 37'b1111111111111101100110111010000110100, 37'b1111111111111010100000101111011001011, 37'b1111111111111111111111000011010111111, 37'b0000000000000000110110110110010010110},
{37'b0000000000000010011101111101011010010, 37'b0000000000000000000001010100000011100, 37'b0000000000000001000011001000000100101, 37'b1111111111111111111111111111110000000, 37'b0000000000000001001110100100000101100, 37'b1111111111111110111011000000011000011, 37'b0000000000000001111000001110000111000, 37'b0000000000000000010101101111000000101, 37'b0000000000000001000101100010100101010, 37'b0000000000000010101110000110000001011, 37'b1111111111111101111001000111111001011, 37'b1111111111111111110101011000000011100, 37'b1111111111111111111011110001011010100, 37'b1111111111111111111011100001000100101, 37'b1111111111111010101110001010011010101, 37'b1111111111111101100111100010100011101, 37'b0000000000000101000010110110100110111, 37'b1111111111111111110001101100110011011, 37'b1111111111111111100101010100101110011, 37'b0000000000000000000000001000010100000, 37'b1111111111111100111101010111011101001, 37'b0000000000000000000100101010011100101, 37'b0000000000000010000000011110100100001, 37'b0000000000000000010011011110110010001, 37'b0000000000000000010010110100010000011, 37'b0000000000000010101101010000110110110, 37'b0000000000000000000000000001000000110, 37'b0000000000000000010011010001010101010, 37'b0000000000000000000000000000000101101, 37'b1111111111111111100111110000011000011, 37'b1111111111111110011001001110001011100, 37'b1111111111111010101011000100111110001, 37'b0000000000000010000111010001100111100, 37'b0000000000000010101111100110011001100, 37'b1111111111111111110001000000010011011, 37'b1111111111111110000111110111010100111, 37'b0000000000000000000000000000101100110, 37'b1111111111111010110000110101111010101, 37'b1111111111111111101000100100010110101, 37'b1111111111111111111110010111100001110, 37'b0000000000000001100100010111111110111, 37'b1111111111111110111101001011101110010, 37'b1111111111111111111111111100010001101, 37'b0000000000000110110001110111000000110, 37'b0000000000000011100101100001011011001, 37'b1111111111111111111100111110001111101, 37'b1111111111111111111111110101010111011, 37'b1111111111111111111111111100010001111, 37'b1111111111111110000100110111111100011, 37'b0000000000000001001011010010100101100, 37'b0000000000000001001001110001110111111, 37'b0000000000000001011001011100000010101, 37'b0000000000000001010000100100011100110, 37'b0000000000000011000110110010101101110, 37'b0000000000000010110011000101001101111, 37'b0000000000000101010001101001111010000, 37'b1111111111111110111000011011001110100, 37'b0000000000000011001001011001010111101, 37'b0000000000000001001110001100010101011, 37'b1111111111111101011001001110100000001, 37'b0000000000000000111000110000001011100, 37'b1111111111111100111001001000010101000, 37'b1111111111111100011110110110110101110, 37'b1111111111111100000000101101101011100},
{37'b0000000000000000000000001010010101101, 37'b0000000000000001110100111101100000110, 37'b1111111111111110011100010111111101010, 37'b0000000000000000000000000010010011110, 37'b1111111111111111100110111001111000010, 37'b1111111111111111101110100011010111111, 37'b1111111111111010101101110100111001111, 37'b1111111111111111111111111100111111011, 37'b0000000000000010000001110000001010100, 37'b0000000000000001111111111010111001100, 37'b0000000000000001111001101110000100011, 37'b1111111111111100110100001010100101100, 37'b1111111111111111010010010101001110101, 37'b0000000000000010010001011010101000011, 37'b1111111111111111111111110110001101110, 37'b0000000000000000000010011100100011100, 37'b1111111111111001010001001101110010111, 37'b1111111111111111111111110101101101100, 37'b0000000000000010111110101111010010010, 37'b0000000000000000100100000110101011011, 37'b0000000000000001111001111010000101010, 37'b1111111111111111000100111111000111011, 37'b0000000000000001111111110100001110110, 37'b0000000000000011001111010101011000110, 37'b1111111111111101001010000110011110100, 37'b1111111111111101110000110010110001100, 37'b1111111111111111111101011000011100001, 37'b1111111111111111010110101000101110011, 37'b0000000000000000100010011011101001101, 37'b0000000000000000000000000100000110111, 37'b1111111111111111111111111101111011000, 37'b0000000000000010100000111001011101000, 37'b1111111111111010000000000110111100111, 37'b0000000000000010111001000001110011101, 37'b0000000000000100000000101110000111010, 37'b0000000000000000111011101011010101110, 37'b0000000000000000111001100101111111100, 37'b1111111111111111001000101111010100011, 37'b0000000000000000111010111110000010101, 37'b1111111111111111001001010110111010000, 37'b1111111111111101111111011001000100111, 37'b1111111111111111100110001110100001001, 37'b0000000000000001010100001101111110011, 37'b0000000000000101100110000101111001010, 37'b1111111111111001001110000111101011110, 37'b1111111111111100011011110010101101001, 37'b0000000000000001100010010111000000011, 37'b1111111111111111001101111000100000101, 37'b0000000000000011100110101100010011100, 37'b1111111111111110000111000110010001010, 37'b1111111111111101010110100000110111001, 37'b1111111111111101110000100001011101000, 37'b1111111111111111111111111110111100110, 37'b0000000000000000111101100100111110110, 37'b1111111111111110101111011110001101111, 37'b1111111111111001010011101000000101111, 37'b1111111111111110110110110010011011111, 37'b1111111111111111111010110001100011011, 37'b0000000000000000010110010010000110110, 37'b1111111111111011000111100011000110101, 37'b0000000000001000111101011110110110100, 37'b1111111111111011101001010100011111001, 37'b0000000000000100010101010110000101111, 37'b0000000000000001001110011100101011101},
{37'b0000000000000000101000000100101001101, 37'b1111111111111110011101110100111011001, 37'b0000000000000101000001101001100101010, 37'b1111111111111101100101001110010110101, 37'b1111111111111100010010110000011111001, 37'b0000000000000000101110000001011010001, 37'b0000000000000010011110011011010001110, 37'b0000000000000010011001111100001011110, 37'b1111111111111110100101001001011000101, 37'b1111111111111110101101110010011111100, 37'b0000000000000000011010111000111101111, 37'b0000000000000001110101010010111000000, 37'b0000000000000001111000010001100011000, 37'b0000000000000000011001101100011010100, 37'b1111111111111110010111011101111011101, 37'b0000000000000001000001110000001010000, 37'b0000000000000011110001000001100010010, 37'b1111111111111111111010010010100001100, 37'b1111111111111101110000110011101001100, 37'b0000000000000000000000000101101001011, 37'b0000000000000000100110000111000111000, 37'b0000000000000000001010011001001101001, 37'b1111111111111101101001111011001010111, 37'b0000000000000000111001110100011111010, 37'b0000000000000110010010111110010100010, 37'b0000000000000000000101001000000110110, 37'b0000000000000001011100011110010000110, 37'b1111111111111001101001111010010000010, 37'b1111111111111111011010110010100011101, 37'b0000000000000000000100110000101100111, 37'b1111111111111110011011100011010011001, 37'b1111111111111101100000011101110000110, 37'b0000000000000011101010101001100010010, 37'b1111111111111111110010011001000001011, 37'b1111111111111111101100101101001110110, 37'b1111111111111101100011110010011000000, 37'b0000000000000001000110111001101001101, 37'b0000000000000010010101100100101111010, 37'b1111111111111111111011000101110000100, 37'b1111111111111111101001110000010001101, 37'b1111111111111110100000011101111011111, 37'b0000000000000001110100111000000011001, 37'b0000000000000000000000000010010001000, 37'b1111111111111010100000100110001100110, 37'b0000000000000010011111010110101101010, 37'b0000000000000011001100010011001100100, 37'b1111111111111111111111111000100001000, 37'b0000000000000000001101000011011001111, 37'b1111111111111100100001110110100110000, 37'b1111111111111111011001101001100010011, 37'b1111111111111111111111111110111110101, 37'b1111111111111101011101011001110101101, 37'b0000000000000000000000000001101011101, 37'b1111111111111110100111100110000010011, 37'b0000000000000000011101010110010111100, 37'b1111111111111001011101100111110001100, 37'b1111111111111111111111111111010101111, 37'b1111111111111111111111100011101100001, 37'b0000000000000010001100111001001011111, 37'b0000000000000100100000010000100011011, 37'b1111111111111010011100001110110011001, 37'b0000000000000100001010010110000100100, 37'b0000000000000000010010111111110100000, 37'b1111111111111111011001110100101111001},
{37'b0000000000000010010011010110111101010, 37'b0000000000001001111011000011101001100, 37'b0000000000000011111101101100100010010, 37'b0000000000000010010010000000011000100, 37'b1111111111111100001011011100011101111, 37'b1111111111111101011101011100100111011, 37'b1111111111101011001101000100100110100, 37'b1111111111111100010110000011110100110, 37'b0000000000000011001110010101001011111, 37'b1111111111111111111111111101000111101, 37'b0000000000000010010110100101001100111, 37'b0000000000000110111001111111101101001, 37'b0000000000000000100011100111010000101, 37'b0000000000000000000010110100001000011, 37'b1111111111111111110111010100000010110, 37'b0000000000000000000000000101100111000, 37'b1111111111111110011111000000011001001, 37'b1111111111111110011000010010001011111, 37'b0000000000000001110101110101100110100, 37'b1111111111111011111110111111001101101, 37'b1111111111111010101011100011001000110, 37'b1111111111111111001011011101111101111, 37'b1111111111111011010101000000011001101, 37'b0000000000000000001111000100000000101, 37'b1111111111101101110010011010101110100, 37'b0000000000000110100001011110101011110, 37'b0000000000000111111010011101101110110, 37'b0000000000000100110101000010100100101, 37'b1111111111110010000011011001010011000, 37'b1111111111111101011111110110110010001, 37'b1111111111111010011111110000110001110, 37'b1111111111111001010000000101100011111, 37'b1111111111101011110011001000101010100, 37'b0000000000000101011010010110001100101, 37'b1111111111111111101001100110110110001, 37'b0000000000000010100011001111000011010, 37'b0000000000000000001100001000011011001, 37'b1111111111110100100010010100111110000, 37'b0000000000000000000000001000110010101, 37'b0000000000000000000000000010101111001, 37'b0000000000000000010000010101100011000, 37'b0000000000001000001001111000111100110, 37'b1111111111111110010111000010010110101, 37'b1111111111111010110101110101110000101, 37'b0000000000000111001011011110010000000, 37'b1111111111111100011100110010100001100, 37'b1111111111111101011001111011011010111, 37'b1111111111111100110111000011101101111, 37'b0000000000000011110100011100101110110, 37'b0000000000000100010000000000000000010, 37'b1111111111111111011101001101010010011, 37'b1111111111111101001101010011101101111, 37'b1111111111111111111110111011000100101, 37'b1111111111111111000110011110100001001, 37'b0000000000000000000000000010100010001, 37'b1111111111111100111110111000100000011, 37'b0000000000000100110110100010001000000, 37'b0000000000001000101011001001001101100, 37'b0000000000000101101100010101110011010, 37'b1111111111111000101110101000111000111, 37'b1111111111100010011000000000011010100, 37'b0000000000000111000101010100111101001, 37'b0000000000000000101111010100100111010, 37'b0000000000000010100010010001101000101},
{37'b1111111111111110000100010100010011010, 37'b0000000000000010101100101100100110000, 37'b0000000000000010100010100110010101010, 37'b1111111111111111111111001100000001111, 37'b1111111111111101000001100101101011001, 37'b1111111111111111010010000101010011110, 37'b1111111111111100111011100100111110101, 37'b1111111111111111100011100000010011100, 37'b0000000000000001001100010101011010000, 37'b1111111111111111011001100100000010101, 37'b1111111111111111110000001011110001100, 37'b1111111111111111101011111101001101110, 37'b1111111111111111111111101001011000111, 37'b1111111111111110100010001001010111010, 37'b1111111111111111110010010110000111001, 37'b1111111111111111001100101000100110101, 37'b0000000000000010100000011111011111001, 37'b1111111111111111111111111111000101100, 37'b1111111111111010110111110010011011110, 37'b0000000000000011101110000110010111001, 37'b0000000000000100110000110110011000111, 37'b0000000000000011010100010011101010010, 37'b1111111111111101011101101011010000000, 37'b1111111111111110111001110111100011010, 37'b1111111111111101001110111000100010000, 37'b1111111111111101101011100110001011100, 37'b0000000000000001110100001110011100111, 37'b0000000000000001110111110001110000110, 37'b0000000000000001110011110001100111001, 37'b0000000000000010111000001110111010100, 37'b0000000000000000010001100001110000001, 37'b0000000000000011000101101011001011101, 37'b1111111111111111101010100100101000001, 37'b0000000000000000000010011110101111101, 37'b0000000000000010011011111110011111110, 37'b0000000000000001000011010110110110001, 37'b1111111111111111011110001101001011111, 37'b1111111111111111111011001001011000001, 37'b0000000000000000000000000011011100000, 37'b1111111111111101101010001101110001001, 37'b1111111111111110001101101010111100000, 37'b1111111111111111000111100001000110101, 37'b1111111111111101001000001011111111111, 37'b0000000000000011100110010010100111110, 37'b0000000000000000000000001001001111000, 37'b1111111111111111111101001010101000111, 37'b1111111111111111010101101100101101001, 37'b1111111111111110110100011011000100100, 37'b1111111111111001100011100011011111000, 37'b1111111111111111101100001000011101110, 37'b1111111111111110001101000110001100010, 37'b1111111111111110110111011100101101001, 37'b1111111111111111001100110111111011111, 37'b0000000000000010000111011010100100000, 37'b0000000000000101011101001101100110000, 37'b0000000000000001011111111110110101011, 37'b1111111111111111111001001100101000010, 37'b1111111111111101010000011010101000011, 37'b1111111111111111110000111100011110000, 37'b0000000000000000000000001010110101011, 37'b0000000000000010100110101111001111111, 37'b1111111111111111110101001010111001101, 37'b0000000000000000010111011111000111010, 37'b0000000000000000000000000000001100000}
};
localparam logic signed [36:0] bias [64] = '{
37'b1111111111111111101100111000000111000,
37'b0000000000000010001100000011111110110,
37'b1111111111111111000000100111101011011,
37'b1111111111111111011110111111110111111,
37'b0000000000000000011011111010110011001,
37'b0000000000000000111011110000100110110,
37'b0000000000000001000101110101110100101,
37'b0000000000000000100110010011111000000,
37'b0000000000000000010111111011100101100,
37'b1111111111111110011000110110100000011,
37'b1111111111111111001101010000101001101,
37'b0000000000000001001101010101011010100,
37'b1111111111111111001011101010100011011,
37'b1111111111111110110101001010110010111,
37'b1111111111111111010011110000010110010,
37'b0000000000000001010101000011111010100,
37'b1111111111111111010101001011101000001,
37'b1111111111111111100010100001101100101,
37'b1111111111111111101111011101110111000,
37'b1111111111111111110001011101110000111,
37'b0000000000000001000000100001100100001,
37'b1111111111111111101101000001011110100,
37'b0000000000000001100011000000001000010,
37'b0000000000000000001010111000000100000,
37'b0000000000000011111111010000111001010,
37'b0000000000000000001000000111000101011,
37'b1111111111111111010101100001011011110,
37'b0000000000000000111000100111000101101,
37'b0000000000000000000110000000101000101,
37'b1111111111111111001000011110101110001,
37'b0000000000000010001100011111010011000,
37'b0000000000000000101111000110100101111,
37'b0000000000000010001100011000111110010,
37'b0000000000000010001010100100001111100,
37'b1111111111111110000000111000000011011,
37'b0000000000000000101000000001111001010,
37'b1111111111111111111101000011100111011,
37'b0000000000000000110111100011011111011,
37'b0000000000000001000101100101101001100,
37'b1111111111111111000010000110110011001,
37'b1111111111111111100010111111001011111,
37'b0000000000000000101111101011001111001,
37'b0000000000000000011100000010111101001,
37'b0000000000000000001111001001011100101,
37'b1111111111111101100000001101011000001,
37'b1111111111111111010100101010000010011,
37'b1111111111111110101010000110111001010,
37'b0000000000000001001011100101010000111,
37'b1111111111111110000111000100101011100,
37'b0000000000000000100001011101101000011,
37'b1111111111111110111110001100010100100,
37'b1111111111111110111001010101010001001,
37'b1111111111111110110010011001011001000,
37'b0000000000000000101000110110110110010,
37'b0000000000000001011100111000101001000,
37'b1111111111111111100100010101001111110,
37'b1111111111111111111010110110100101100,
37'b0000000000000000100001110110010111100,
37'b0000000000000000011001110111111000110,
37'b0000000000000000001101110000001011010,
37'b0000000000000000010000110011111011010,
37'b0000000000000001001111101010001001100,
37'b1111111111111101101101011001001111111,
37'b1111111111111111010011000110100010101
};
endpackage