// Package with weights and biases for pre-sigmoid dense latency layer
`ifndef DENSE_LAYER_1_PKG
    `define DENSE_LAYER_1_PKG dense_1_gen
`endif

`ifndef DENSE_LAYER_2_PKG
    `define DENSE_LAYER_2_PKG dense_2_gen
`endif

`ifndef DENSE_LAYER_3_PKG
    `define DENSE_LAYER_3_PKG dense_3_gen
`endif

`ifndef DENSE_LAYER_4_PKG
    `define DENSE_LAYER_4_PKG dense_4_gen
`endif