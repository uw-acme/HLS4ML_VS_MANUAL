// Width: 14
// NFRAC: 7
package dense_1_14_7;

localparam logic signed [13:0] weights [16][64] = '{ 
{14'b00000000100000, 14'b11111110101100, 14'b11111111101000, 14'b11111111100011, 14'b11111111001100, 14'b00000000001110, 14'b11111101111011, 14'b00000000000000, 14'b00000000000111, 14'b00000000100001, 14'b00000000000000, 14'b11111111001100, 14'b11111111111111, 14'b00000000011010, 14'b00000000000100, 14'b11111111011110, 14'b00000000011101, 14'b00000000000111, 14'b00000000000000, 14'b11111111111111, 14'b00000000110000, 14'b11111111010101, 14'b11111111111101, 14'b00000000111100, 14'b11111111010110, 14'b11111110101000, 14'b11111111011100, 14'b11111111100111, 14'b11111111110010, 14'b11111111111111, 14'b00000000000100, 14'b00000000011111, 14'b00000000011001, 14'b11111111111110, 14'b00000000000000, 14'b00000000100111, 14'b11111111111101, 14'b11111111011111, 14'b00000000000011, 14'b00000000011000, 14'b11111111111110, 14'b00000000100011, 14'b11111111011101, 14'b00000001110110, 14'b11111111111111, 14'b00000000111001, 14'b00000000000000, 14'b00000000010111, 14'b00000000011001, 14'b11111111111100, 14'b00000000000000, 14'b00000000010100, 14'b00000000011011, 14'b00000000001001, 14'b11111111110001, 14'b11111111011000, 14'b00000001000100, 14'b11111111000000, 14'b00000000111011, 14'b11111111010010, 14'b00000001100101, 14'b11111111111111, 14'b00000000000001, 14'b00000000001010}, 
{14'b00000000000000, 14'b11111111010110, 14'b11111111101111, 14'b11111111011100, 14'b11111111010111, 14'b00000000001101, 14'b11111110011111, 14'b11111111111111, 14'b11111111100010, 14'b00000000010110, 14'b00000000000000, 14'b11111111110100, 14'b00000000011001, 14'b00000000000000, 14'b11111111111111, 14'b00000000011010, 14'b11111111111111, 14'b00000000000000, 14'b11111111101000, 14'b11111111011111, 14'b00000000111000, 14'b11111111110101, 14'b00000000000110, 14'b00000001011001, 14'b00000000100000, 14'b11111111100010, 14'b11111111100010, 14'b11111111111111, 14'b11111111110011, 14'b11111111001100, 14'b11111111111000, 14'b00000000111010, 14'b00000000100011, 14'b00000001000110, 14'b00000001010000, 14'b00000000000110, 14'b11111111110000, 14'b11111111001000, 14'b00000000000111, 14'b00000000011000, 14'b00000000000010, 14'b00000000011010, 14'b11111111100100, 14'b00000000100000, 14'b00000000010110, 14'b00000000000110, 14'b11111111010100, 14'b00000000001010, 14'b00000000100001, 14'b00000000000011, 14'b00000000000011, 14'b00000010010100, 14'b11111111110110, 14'b11111111110011, 14'b11111111111001, 14'b11111111111111, 14'b00000000100000, 14'b11111111010000, 14'b00000001111110, 14'b00000000000000, 14'b00000001000010, 14'b00000000011110, 14'b00000001101001, 14'b00000000010010}, 
{14'b11111111111111, 14'b00000000000000, 14'b11111111110101, 14'b11111111101001, 14'b11111111101000, 14'b00000000000101, 14'b00000010111101, 14'b11111111111111, 14'b11111101011101, 14'b11111111111111, 14'b11111111111111, 14'b11111111111101, 14'b11111111100010, 14'b00000000000000, 14'b11111111111110, 14'b00000000010101, 14'b00000001110011, 14'b11111111111111, 14'b00000000001001, 14'b00000000000000, 14'b00000000110100, 14'b11111110100011, 14'b00000001001001, 14'b11111110100100, 14'b00000001111001, 14'b11111111010011, 14'b11111111100000, 14'b11111110100100, 14'b00000010100011, 14'b00000000100011, 14'b00000000000001, 14'b00000001000010, 14'b00000010000010, 14'b11111101100111, 14'b11111111110011, 14'b00000000000100, 14'b11111111100010, 14'b00000001110010, 14'b11111111111010, 14'b00000000101000, 14'b00000000101010, 14'b00000000101111, 14'b11111111111111, 14'b11111111111111, 14'b11111111111101, 14'b00000000010100, 14'b11111111011100, 14'b11111111101010, 14'b11111111111101, 14'b00000000110010, 14'b11111111101001, 14'b00000000010011, 14'b11111111111111, 14'b00000000010001, 14'b11111111101001, 14'b11111111111111, 14'b11111111011000, 14'b11111110101010, 14'b11111111111111, 14'b00000000000000, 14'b00000011000101, 14'b00000000000001, 14'b11111111111111, 14'b11111111011000}, 
{14'b11111111000101, 14'b11111111010000, 14'b11111110100111, 14'b00000000100111, 14'b11111111010111, 14'b11111101010011, 14'b11111111110001, 14'b11111111011000, 14'b00000000011100, 14'b11111111111111, 14'b00000010100001, 14'b11111111110010, 14'b11111110011011, 14'b00000001001010, 14'b00000000000011, 14'b11111111111111, 14'b11111111000111, 14'b11111111111111, 14'b00000000000000, 14'b11111111100011, 14'b11111101101100, 14'b11111111110001, 14'b11111110100110, 14'b00000000011001, 14'b11111111001110, 14'b11111110001010, 14'b00000000101000, 14'b00000001011110, 14'b00000010100101, 14'b11111111000101, 14'b11111110110101, 14'b00000000001001, 14'b00000001000000, 14'b11111110010100, 14'b11111111010111, 14'b00000000000000, 14'b11111110100011, 14'b00000000011111, 14'b11111111000111, 14'b00000000001111, 14'b00000000111010, 14'b00000000010100, 14'b00000000000000, 14'b00000000000010, 14'b00000001000110, 14'b11111111100110, 14'b11111111111111, 14'b11111111010011, 14'b11111111111111, 14'b11111111110011, 14'b11111110110001, 14'b00000000001011, 14'b11111111111111, 14'b00000000011011, 14'b00000000101000, 14'b00000001010010, 14'b11111110000100, 14'b11111110001001, 14'b11111110100101, 14'b00000001101110, 14'b00000011011111, 14'b11111110001100, 14'b11111111111001, 14'b00000000110111}, 
{14'b00000000101011, 14'b11111110110000, 14'b11111111011110, 14'b11111111111111, 14'b11111111101100, 14'b00000000101011, 14'b00000000011000, 14'b11111111111111, 14'b11111110110011, 14'b11111111100001, 14'b11111111010000, 14'b00000000000110, 14'b00000000000000, 14'b00000000000000, 14'b11111111111010, 14'b00000000101101, 14'b00000000010001, 14'b11111111001101, 14'b00000000000011, 14'b00000000000001, 14'b00000000011010, 14'b11111111110000, 14'b00000000001001, 14'b11111111111101, 14'b00000010001000, 14'b11111111101000, 14'b11111111011100, 14'b11111111001100, 14'b00000000000000, 14'b00000000010101, 14'b00000000001110, 14'b00000000100011, 14'b11111111111110, 14'b00000000001001, 14'b00000000010000, 14'b11111111111111, 14'b00000000000000, 14'b00000001110000, 14'b11111111011011, 14'b11111111110110, 14'b00000000110111, 14'b00000000011111, 14'b11111111000001, 14'b00000000000000, 14'b11111101110111, 14'b11111111111111, 14'b11111111110000, 14'b00000000000001, 14'b11111111111111, 14'b11111111111100, 14'b11111111111111, 14'b00000000011000, 14'b11111111111111, 14'b00000000101000, 14'b11111111100111, 14'b11111110100001, 14'b11111111000100, 14'b11111110111110, 14'b11111110110001, 14'b00000001011111, 14'b00000010101111, 14'b00000001100101, 14'b00000000001111, 14'b11111111111111}, 
{14'b11111111000110, 14'b11111110101111, 14'b00000000000000, 14'b00000000100111, 14'b00000000100100, 14'b11111111100100, 14'b00000001001010, 14'b11111111111111, 14'b00000000011111, 14'b11111111111111, 14'b11111111111110, 14'b11111111110110, 14'b11111111101001, 14'b00000001001010, 14'b11111111110100, 14'b00000000000000, 14'b11111110110000, 14'b11111111010010, 14'b00000000000000, 14'b11111111111111, 14'b11111111111001, 14'b11111111010111, 14'b11111111010111, 14'b00000000111011, 14'b11111111010111, 14'b11111111111111, 14'b00000000100000, 14'b11111111110110, 14'b11111110001000, 14'b11111111111111, 14'b11111111110111, 14'b11111111111110, 14'b11111111111110, 14'b00000000000101, 14'b00000000010000, 14'b00000000101100, 14'b00000000000001, 14'b11111111110011, 14'b11111111011110, 14'b11111111111111, 14'b11111111101010, 14'b11111110111100, 14'b00000000110011, 14'b00000000000001, 14'b00000001001101, 14'b00000000000000, 14'b11111111111111, 14'b00000000001100, 14'b11111111001010, 14'b00000000011101, 14'b00000000000000, 14'b11111111110011, 14'b11111111010001, 14'b00000000110001, 14'b11111111111111, 14'b00000000101100, 14'b00000000011011, 14'b00000000011010, 14'b11111111111101, 14'b11111111111110, 14'b11111110011000, 14'b11111111101111, 14'b11111111111000, 14'b11111111111111}, 
{14'b11111111011011, 14'b11111111010101, 14'b11111111001000, 14'b11111111110111, 14'b11111111101110, 14'b00000000001101, 14'b11111110100110, 14'b11111111101100, 14'b11111111100011, 14'b11111111111111, 14'b11111111011011, 14'b00000000101100, 14'b00000000000100, 14'b00000000010001, 14'b00000000100111, 14'b00000000000000, 14'b00000001100110, 14'b00000000001011, 14'b00000000011111, 14'b00000000100010, 14'b11111111101011, 14'b00000000101110, 14'b11111111100000, 14'b11111110111111, 14'b00000000010110, 14'b00000001000010, 14'b11111111111111, 14'b00000000000110, 14'b11111110000110, 14'b00000000100100, 14'b00000000100010, 14'b11111111010000, 14'b00000000111100, 14'b00000001010101, 14'b00000000000000, 14'b00000000101011, 14'b11111111111111, 14'b00000000100100, 14'b00000000011001, 14'b00000000000000, 14'b11111111110000, 14'b11111111010001, 14'b00000000010010, 14'b00000000111101, 14'b00000001000010, 14'b11111111101010, 14'b11111111110101, 14'b11111111100111, 14'b11111111101110, 14'b00000000001111, 14'b00000000000000, 14'b00000000000100, 14'b00000000000000, 14'b00000000010111, 14'b11111111101001, 14'b00000001100010, 14'b00000000101101, 14'b11111111111100, 14'b00000000110001, 14'b00000000011011, 14'b11111100101111, 14'b11111110110110, 14'b11111111101001, 14'b11111111111110}, 
{14'b00000000000000, 14'b00000000011110, 14'b11111111111111, 14'b11111111111111, 14'b11111111010110, 14'b11111111111100, 14'b11111111011111, 14'b00000000000000, 14'b00000000000011, 14'b00000000110001, 14'b00000000000001, 14'b11111111001111, 14'b11111111110111, 14'b00000000000000, 14'b11111111111001, 14'b11111111000110, 14'b11111110010011, 14'b11111111111111, 14'b11111110110010, 14'b11111111000110, 14'b11111111001110, 14'b00000000101100, 14'b00000000000110, 14'b11111111101101, 14'b11111111001000, 14'b00000000010011, 14'b00000000000000, 14'b00000000111111, 14'b00000001100111, 14'b11111111111010, 14'b00000000000000, 14'b00000000011101, 14'b11111110101000, 14'b11111111010000, 14'b00000000000111, 14'b00000000001011, 14'b11111111011100, 14'b00000000011110, 14'b00000000010000, 14'b11111111101100, 14'b11111111001010, 14'b11111111111011, 14'b00000000000100, 14'b11111111101010, 14'b00000000000111, 14'b00000000011101, 14'b11111111110000, 14'b00000000000011, 14'b00000000000000, 14'b11111111100100, 14'b11111111001110, 14'b00000000110101, 14'b00000000010000, 14'b11111111101001, 14'b00000000010000, 14'b11111111111000, 14'b11111111000011, 14'b11111111101110, 14'b11111111111001, 14'b11111111110111, 14'b00000001101010, 14'b00000000011000, 14'b11111111111001, 14'b11111111111111}, 
{14'b00000000000001, 14'b00000001001011, 14'b11111110110101, 14'b11111111100010, 14'b00000000101001, 14'b11111111100101, 14'b00000010011011, 14'b11111111011011, 14'b11111111111111, 14'b00000000100101, 14'b00000000100000, 14'b11111111111111, 14'b11111111111001, 14'b11111111000010, 14'b00000000100100, 14'b00000000010100, 14'b11111111100111, 14'b11111111111111, 14'b00000000000000, 14'b00000000000000, 14'b00000000100001, 14'b11111111000101, 14'b00000000110010, 14'b00000001001110, 14'b11111111110100, 14'b11111111111111, 14'b11111111111101, 14'b11111111111111, 14'b00000001011110, 14'b00000000000000, 14'b11111111011101, 14'b00000000000000, 14'b00000000110001, 14'b11111110011000, 14'b11111110111010, 14'b00000000011001, 14'b00000000010001, 14'b11111110110110, 14'b11111111100111, 14'b11111111100100, 14'b00000000110011, 14'b00000000110010, 14'b00000000000000, 14'b11111111011101, 14'b00000000000000, 14'b00000000110010, 14'b11111111111000, 14'b11111111111111, 14'b00000000000001, 14'b00000000011111, 14'b11111111111000, 14'b11111111100111, 14'b00000000101100, 14'b11111111100100, 14'b00000000100011, 14'b00000001001010, 14'b00000000000101, 14'b00000000100001, 14'b11111111001100, 14'b11111111010001, 14'b00000001101010, 14'b11111111101111, 14'b00000000000101, 14'b11111111110100}, 
{14'b00000000000010, 14'b11111111000110, 14'b00000000101111, 14'b11111111011011, 14'b11111111111111, 14'b00000000011011, 14'b11111110110101, 14'b00000000011000, 14'b00000000111110, 14'b00000000010011, 14'b00000000101110, 14'b00000000101001, 14'b11111111011000, 14'b11111111110110, 14'b11111111111001, 14'b00000000000000, 14'b11111110000101, 14'b00000000101001, 14'b11111111111011, 14'b00000000000011, 14'b11111111010010, 14'b00000000001000, 14'b00000000010011, 14'b11111111111111, 14'b11111111000101, 14'b11111111111001, 14'b11111111110101, 14'b00000010011111, 14'b11111110101011, 14'b00000000001000, 14'b00000000001100, 14'b11111111111000, 14'b11111111100011, 14'b00000000001110, 14'b11111111110101, 14'b11111111101110, 14'b11111111101001, 14'b11111111100101, 14'b11111111111101, 14'b11111111011001, 14'b00000000101001, 14'b00000000001111, 14'b00000000111111, 14'b00000000001011, 14'b00000000000100, 14'b11111111011010, 14'b00000000000000, 14'b11111111111111, 14'b11111111111111, 14'b00000000011000, 14'b00000000010110, 14'b00000000100101, 14'b11111111111111, 14'b11111111011010, 14'b00000000000001, 14'b00000000000000, 14'b00000000101001, 14'b11111111100110, 14'b11111110111001, 14'b00000001000111, 14'b11111111011010, 14'b00000010010100, 14'b11111111111101, 14'b11111111010010}, 
{14'b11111110110110, 14'b11111111111111, 14'b11111111001011, 14'b00000000011101, 14'b00000000100001, 14'b11111111110010, 14'b00000001000010, 14'b11111111101010, 14'b11111111000010, 14'b11111111010001, 14'b11111111011111, 14'b11111111000011, 14'b11111111100010, 14'b00000000011001, 14'b00000000000000, 14'b00000000000000, 14'b00000001101011, 14'b11111111111010, 14'b11111111111111, 14'b00000000110100, 14'b00000000100101, 14'b11111110110101, 14'b11111111001111, 14'b00000000011000, 14'b11111111001000, 14'b11111111111101, 14'b11111111011110, 14'b11111111010101, 14'b11111111001000, 14'b00000000100110, 14'b00000000011101, 14'b11111111101100, 14'b11111111110110, 14'b11111110000011, 14'b11111111101001, 14'b00000000000110, 14'b11111111101111, 14'b11111111011010, 14'b11111111111111, 14'b00000000001111, 14'b11111111110000, 14'b11111111111111, 14'b11111111111011, 14'b11111110101010, 14'b00000000000000, 14'b00000000000000, 14'b00000000101011, 14'b11111111110000, 14'b00000000110110, 14'b11111111100111, 14'b00000000100100, 14'b11111111111111, 14'b00000000011100, 14'b11111111001101, 14'b11111111111111, 14'b00000001000001, 14'b00000000101000, 14'b00000000100101, 14'b00000000000011, 14'b11111111001100, 14'b11111111011001, 14'b11111110101000, 14'b11111111111111, 14'b00000000001101}, 
{14'b00000000100111, 14'b00000000000000, 14'b00000000010000, 14'b11111111111111, 14'b00000000010011, 14'b11111111101110, 14'b00000000011110, 14'b00000000000101, 14'b00000000010001, 14'b00000000101011, 14'b11111111011110, 14'b11111111111101, 14'b11111111111110, 14'b11111111111110, 14'b11111110101011, 14'b11111111011001, 14'b00000001010000, 14'b11111111111100, 14'b11111111111001, 14'b00000000000000, 14'b11111111001111, 14'b00000000000001, 14'b00000000100000, 14'b00000000000100, 14'b00000000000100, 14'b00000000101011, 14'b00000000000000, 14'b00000000000100, 14'b00000000000000, 14'b11111111111001, 14'b11111111100110, 14'b11111110101010, 14'b00000000100001, 14'b00000000101011, 14'b11111111111100, 14'b11111111100001, 14'b00000000000000, 14'b11111110101100, 14'b11111111111010, 14'b11111111111111, 14'b00000000011001, 14'b11111111101111, 14'b11111111111111, 14'b00000001101100, 14'b00000000111001, 14'b11111111111111, 14'b11111111111111, 14'b11111111111111, 14'b11111111100001, 14'b00000000010010, 14'b00000000010010, 14'b00000000010110, 14'b00000000010100, 14'b00000000110001, 14'b00000000101100, 14'b00000001010100, 14'b11111111101110, 14'b00000000110010, 14'b00000000010011, 14'b11111111010110, 14'b00000000001110, 14'b11111111001110, 14'b11111111000111, 14'b11111111000000}, 
{14'b00000000000000, 14'b00000000011101, 14'b11111111100111, 14'b00000000000000, 14'b11111111111001, 14'b11111111111011, 14'b11111110101011, 14'b11111111111111, 14'b00000000100000, 14'b00000000011111, 14'b00000000011110, 14'b11111111001101, 14'b11111111110100, 14'b00000000100100, 14'b11111111111111, 14'b00000000000000, 14'b11111110010100, 14'b11111111111111, 14'b00000000101111, 14'b00000000001001, 14'b00000000011110, 14'b11111111110001, 14'b00000000011111, 14'b00000000110011, 14'b11111111010010, 14'b11111111011100, 14'b11111111111111, 14'b11111111110101, 14'b00000000001000, 14'b00000000000000, 14'b11111111111111, 14'b00000000101000, 14'b11111110100000, 14'b00000000101110, 14'b00000001000000, 14'b00000000001110, 14'b00000000001110, 14'b11111111110010, 14'b00000000001110, 14'b11111111110010, 14'b11111111011111, 14'b11111111111001, 14'b00000000010101, 14'b00000001011001, 14'b11111110010011, 14'b11111111000110, 14'b00000000011000, 14'b11111111110011, 14'b00000000111001, 14'b11111111100001, 14'b11111111010101, 14'b11111111011100, 14'b11111111111111, 14'b00000000001111, 14'b11111111101011, 14'b11111110010100, 14'b11111111101101, 14'b11111111111110, 14'b00000000000101, 14'b11111110110001, 14'b00000010001111, 14'b11111110111010, 14'b00000001000101, 14'b00000000010011}, 
{14'b00000000001010, 14'b11111111100111, 14'b00000001010000, 14'b11111111011001, 14'b11111111000100, 14'b00000000001011, 14'b00000000100111, 14'b00000000100110, 14'b11111111101001, 14'b11111111101011, 14'b00000000000110, 14'b00000000011101, 14'b00000000011110, 14'b00000000000110, 14'b11111111100101, 14'b00000000010000, 14'b00000000111100, 14'b11111111111110, 14'b11111111011100, 14'b00000000000000, 14'b00000000001001, 14'b00000000000010, 14'b11111111011010, 14'b00000000001110, 14'b00000001100100, 14'b00000000000001, 14'b00000000010111, 14'b11111110011010, 14'b11111111110110, 14'b00000000000001, 14'b11111111100110, 14'b11111111011000, 14'b00000000111010, 14'b11111111111100, 14'b11111111111011, 14'b11111111011000, 14'b00000000010001, 14'b00000000100101, 14'b11111111111110, 14'b11111111111010, 14'b11111111101000, 14'b00000000011101, 14'b00000000000000, 14'b11111110101000, 14'b00000000100111, 14'b00000000110011, 14'b11111111111111, 14'b00000000000011, 14'b11111111001000, 14'b11111111110110, 14'b11111111111111, 14'b11111111010111, 14'b00000000000000, 14'b11111111101001, 14'b00000000000111, 14'b11111110010111, 14'b11111111111111, 14'b11111111111111, 14'b00000000100011, 14'b00000001001000, 14'b11111110100111, 14'b00000001000010, 14'b00000000000100, 14'b11111111110110}, 
{14'b00000000100100, 14'b00000010011110, 14'b00000000111111, 14'b00000000100100, 14'b11111111000010, 14'b11111111010111, 14'b11111010110011, 14'b11111111000101, 14'b00000000110011, 14'b11111111111111, 14'b00000000100101, 14'b00000001101110, 14'b00000000001000, 14'b00000000000000, 14'b11111111111101, 14'b00000000000000, 14'b11111111100111, 14'b11111111100110, 14'b00000000011101, 14'b11111110111111, 14'b11111110101010, 14'b11111111110010, 14'b11111110110101, 14'b00000000000011, 14'b11111011011100, 14'b00000001101000, 14'b00000001111110, 14'b00000001001101, 14'b11111100100000, 14'b11111111010111, 14'b11111110100111, 14'b11111110010100, 14'b11111010111100, 14'b00000001010110, 14'b11111111111010, 14'b00000000101000, 14'b00000000000011, 14'b11111101001000, 14'b00000000000000, 14'b00000000000000, 14'b00000000000100, 14'b00000010000010, 14'b11111111100101, 14'b11111110101101, 14'b00000001110010, 14'b11111111000111, 14'b11111111010110, 14'b11111111001101, 14'b00000000111101, 14'b00000001000100, 14'b11111111110111, 14'b11111111010011, 14'b11111111111111, 14'b11111111110001, 14'b00000000000000, 14'b11111111001111, 14'b00000001001101, 14'b00000010001010, 14'b00000001011011, 14'b11111110001011, 14'b11111000100110, 14'b00000001110001, 14'b00000000001011, 14'b00000000101000}, 
{14'b11111111100001, 14'b00000000101011, 14'b00000000101000, 14'b11111111111111, 14'b11111111010000, 14'b11111111110100, 14'b11111111001110, 14'b11111111111000, 14'b00000000010011, 14'b11111111110110, 14'b11111111111100, 14'b11111111111010, 14'b11111111111111, 14'b11111111101000, 14'b11111111111100, 14'b11111111110011, 14'b00000000101000, 14'b11111111111111, 14'b11111110101101, 14'b00000000111011, 14'b00000001001100, 14'b00000000110101, 14'b11111111010111, 14'b11111111101110, 14'b11111111010011, 14'b11111111011010, 14'b00000000011101, 14'b00000000011101, 14'b00000000011100, 14'b00000000101110, 14'b00000000000100, 14'b00000000110001, 14'b11111111111010, 14'b00000000000000, 14'b00000000100110, 14'b00000000010000, 14'b11111111110111, 14'b11111111111110, 14'b00000000000000, 14'b11111111011010, 14'b11111111100011, 14'b11111111110001, 14'b11111111010010, 14'b00000000111001, 14'b00000000000000, 14'b11111111111111, 14'b11111111110101, 14'b11111111101101, 14'b11111110011000, 14'b11111111111011, 14'b11111111100011, 14'b11111111101101, 14'b11111111110011, 14'b00000000100001, 14'b00000001010111, 14'b00000000010111, 14'b11111111111110, 14'b11111111010100, 14'b11111111111100, 14'b00000000000000, 14'b00000000101001, 14'b11111111111101, 14'b00000000000101, 14'b00000000000000}
};

localparam logic signed [13:0] bias [64] = '{
14'b11111111111011,  // -0.037350185215473175
14'b00000000100011,  // 0.27355897426605225
14'b11111111110000,  // -0.12378914654254913
14'b11111111110111,  // -0.064457006752491
14'b00000000000110,  // 0.05452875792980194
14'b00000000001110,  // 0.11671770364046097
14'b00000000010001,  // 0.13640816509723663
14'b00000000001001,  // 0.07482525706291199
14'b00000000000101,  // 0.04674031585454941
14'b11111111100110,  // -0.20146161317825317
14'b11111111110011,  // -0.09910125285387039
14'b00000000010011,  // 0.15104414522647858
14'b11111111110010,  // -0.10221704095602036
14'b11111111101101,  // -0.1461549550294876
14'b11111111110100,  // -0.08641516417264938
14'b00000000010101,  // 0.16613510251045227
14'b11111111110101,  // -0.0836295336484909
14'b11111111111000,  // -0.05756539851427078
14'b11111111111011,  // -0.03229188174009323
14'b11111111111100,  // -0.028388574719429016
14'b00000000010000,  // 0.1260243058204651
14'b11111111111011,  // -0.037064336240291595
14'b00000000011000,  // 0.19336333870887756
14'b00000000000010,  // 0.02124214917421341
14'b00000000111111,  // 0.4985624849796295
14'b00000000000010,  // 0.0158411655575037
14'b11111111110101,  // -0.08296407759189606
14'b00000000001110,  // 0.11056788265705109
14'b00000000000001,  // 0.01173810102045536
14'b11111111110010,  // -0.10843746364116669
14'b00000000100011,  // 0.27439257502555847
14'b00000000001011,  // 0.09199801832437515
14'b00000000100011,  // 0.27419957518577576
14'b00000000100010,  // 0.27063727378845215
14'b11111111100000,  // -0.24828937649726868
14'b00000000001010,  // 0.07818280160427094
14'b11111111111111,  // -0.005749030504375696
14'b00000000001101,  // 0.10850494354963303
14'b00000000010001,  // 0.13591453433036804
14'b11111111110000,  // -0.12088628858327866
14'b11111111111000,  // -0.05666546896100044
14'b00000000001011,  // 0.09311636537313461
14'b00000000000111,  // 0.05477767437696457
14'b00000000000011,  // 0.029585206881165504
14'b11111111011000,  // -0.31209176778793335
14'b11111111110101,  // -0.08465463668107986
14'b11111111101010,  // -0.16775836050510406
14'b00000000010010,  // 0.14762157201766968
14'b11111111100001,  // -0.23618532717227936
14'b00000000001000,  // 0.06535740196704865
14'b11111111101111,  // -0.12853026390075684
14'b11111111101110,  // -0.13802281022071838
14'b11111111101100,  // -0.15156887471675873
14'b00000000001010,  // 0.07979883998632431
14'b00000000010111,  // 0.18141601979732513
14'b11111111111001,  // -0.054039113223552704
14'b11111111111110,  // -0.010052933357656002
14'b00000000001000,  // 0.06611225008964539
14'b00000000000110,  // 0.05053366720676422
14'b00000000000011,  // 0.026860840618610382
14'b00000000000100,  // 0.03283466026186943
14'b00000000010011,  // 0.15558314323425293
14'b11111111011011,  // -0.2863388657569885
14'b11111111110100   // -0.08769102394580841
};
endpackage