//Width: 4
//Int: 2
package dense_4_gen;

localparam logic signed [3:0] weights [32][5] = '{
{4'b1111, 4'b0001, 4'b1111, 4'b0000, 4'b1111},
{4'b1110, 4'b1111, 4'b0010, 4'b1111, 4'b0000},
{4'b0001, 4'b0001, 4'b1111, 4'b1110, 4'b1111},
{4'b1110, 4'b1111, 4'b1111, 4'b0001, 4'b0001},
{4'b0000, 4'b0001, 4'b0001, 4'b1111, 4'b1100},
{4'b0001, 4'b1110, 4'b0001, 4'b1111, 4'b1111},
{4'b1110, 4'b0000, 4'b1111, 4'b0001, 4'b0000},
{4'b1111, 4'b0001, 4'b1110, 4'b0001, 4'b0001},
{4'b0001, 4'b1111, 4'b0000, 4'b1110, 4'b1111},
{4'b1111, 4'b1111, 4'b0001, 4'b0010, 4'b0000},
{4'b1111, 4'b1111, 4'b0000, 4'b0010, 4'b1111},
{4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b0000},
{4'b0000, 4'b0001, 4'b0000, 4'b1111, 4'b1110},
{4'b0001, 4'b0000, 4'b0010, 4'b1111, 4'b1110},
{4'b0000, 4'b1111, 4'b1111, 4'b1111, 4'b0010},
{4'b1110, 4'b1111, 4'b1111, 4'b0010, 4'b0000},
{4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b1111},
{4'b0001, 4'b1111, 4'b1110, 4'b1111, 4'b0000},
{4'b0001, 4'b0000, 4'b1111, 4'b0000, 4'b1110},
{4'b0001, 4'b1111, 4'b1111, 4'b0001, 4'b0000},
{4'b0000, 4'b1111, 4'b0001, 4'b1110, 4'b1111},
{4'b0000, 4'b0000, 4'b0010, 4'b1110, 4'b1110},
{4'b1111, 4'b0000, 4'b0001, 4'b1111, 4'b0010},
{4'b1111, 4'b0001, 4'b0001, 4'b0000, 4'b1110},
{4'b1111, 4'b0001, 4'b1111, 4'b0000, 4'b0010},
{4'b0000, 4'b0001, 4'b0000, 4'b1101, 4'b0010},
{4'b1110, 4'b1111, 4'b0001, 4'b0001, 4'b0001},
{4'b0000, 4'b0001, 4'b1111, 4'b1111, 4'b0000},
{4'b1111, 4'b0001, 4'b1110, 4'b0001, 4'b1111},
{4'b1111, 4'b0001, 4'b1111, 4'b1110, 4'b0010},
{4'b0010, 4'b0000, 4'b0001, 4'b1110, 4'b1111},
{4'b1111, 4'b1110, 4'b0001, 4'b0000, 4'b0001}
};
localparam logic signed [3:0] bias [5] = '{
4'b1111,
4'b1111,
4'b1111,
4'b0000,
4'b0001
};
endpackage